VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO audiodac_drv
  CLASS BLOCK ;
  FOREIGN audiodac_drv ;
  ORIGIN -0.105 0.000 ;
  SIZE 73.715 BY 141.930 ;
  PIN in_p
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 3.265 62.940 3.595 63.110 ;
        RECT 4.225 62.940 4.555 63.110 ;
        RECT 5.175 62.940 5.505 63.110 ;
        RECT 6.135 62.940 6.465 63.110 ;
        RECT 7.095 62.940 7.425 63.110 ;
        RECT 2.785 60.390 3.115 60.560 ;
        RECT 3.745 60.390 4.075 60.560 ;
        RECT 4.705 60.390 5.035 60.560 ;
        RECT 5.655 60.390 5.985 60.560 ;
        RECT 6.615 60.390 6.945 60.560 ;
      LAYER mcon ;
        RECT 3.345 62.940 3.515 63.110 ;
        RECT 4.305 62.940 4.475 63.110 ;
        RECT 5.255 62.940 5.425 63.110 ;
        RECT 6.215 62.940 6.385 63.110 ;
        RECT 7.175 62.940 7.345 63.110 ;
        RECT 2.865 60.390 3.035 60.560 ;
        RECT 3.825 60.390 3.995 60.560 ;
        RECT 4.785 60.390 4.955 60.560 ;
        RECT 5.735 60.390 5.905 60.560 ;
        RECT 6.695 60.390 6.865 60.560 ;
      LAYER met1 ;
        RECT 1.965 62.905 7.615 63.145 ;
        RECT 1.965 62.045 2.215 62.905 ;
        RECT 1.855 61.645 2.325 62.045 ;
        RECT 1.965 61.515 2.215 61.645 ;
        RECT 1.975 60.595 2.215 61.515 ;
        RECT 1.975 60.355 7.615 60.595 ;
      LAYER via ;
        RECT 1.905 61.645 2.275 62.045 ;
      LAYER met2 ;
        RECT 1.905 61.595 2.275 62.095 ;
      LAYER via2 ;
        RECT 1.905 61.645 2.275 62.045 ;
      LAYER met3 ;
        RECT 1.855 62.045 2.325 62.070 ;
        RECT 0.455 61.645 14.155 62.045 ;
        RECT 1.855 61.620 2.325 61.645 ;
    END
  END in_p
  PIN in_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 9.195 62.940 9.525 63.110 ;
        RECT 10.155 62.940 10.485 63.110 ;
        RECT 11.105 62.940 11.435 63.110 ;
        RECT 12.065 62.940 12.395 63.110 ;
        RECT 13.025 62.940 13.355 63.110 ;
        RECT 8.715 60.390 9.045 60.560 ;
        RECT 9.675 60.390 10.005 60.560 ;
        RECT 10.635 60.390 10.965 60.560 ;
        RECT 11.585 60.390 11.915 60.560 ;
        RECT 12.545 60.390 12.875 60.560 ;
      LAYER mcon ;
        RECT 9.275 62.940 9.445 63.110 ;
        RECT 10.235 62.940 10.405 63.110 ;
        RECT 11.185 62.940 11.355 63.110 ;
        RECT 12.145 62.940 12.315 63.110 ;
        RECT 13.105 62.940 13.275 63.110 ;
        RECT 8.795 60.390 8.965 60.560 ;
        RECT 9.755 60.390 9.925 60.560 ;
        RECT 10.715 60.390 10.885 60.560 ;
        RECT 11.665 60.390 11.835 60.560 ;
        RECT 12.625 60.390 12.795 60.560 ;
      LAYER met1 ;
        RECT 8.515 62.945 14.155 63.145 ;
        RECT 8.515 62.905 14.275 62.945 ;
        RECT 13.805 62.545 14.275 62.905 ;
        RECT 13.915 60.595 14.155 62.545 ;
        RECT 8.515 60.355 14.155 60.595 ;
      LAYER via ;
        RECT 13.855 62.545 14.225 62.945 ;
      LAYER met2 ;
        RECT 13.855 62.495 14.225 62.995 ;
      LAYER via2 ;
        RECT 13.855 62.545 14.225 62.945 ;
      LAYER met3 ;
        RECT 13.805 62.945 14.275 62.970 ;
        RECT 0.455 62.545 14.275 62.945 ;
        RECT 13.805 62.520 14.275 62.545 ;
    END
  END in_n
  PIN out_p
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 435.000000 ;
    PORT
      LAYER li1 ;
        RECT 26.035 59.115 26.205 69.155 ;
        RECT 27.615 59.115 27.785 69.155 ;
        RECT 29.195 59.115 29.365 69.155 ;
        RECT 30.775 59.115 30.945 69.155 ;
        RECT 32.355 59.115 32.525 69.155 ;
        RECT 35.975 59.115 36.145 69.155 ;
        RECT 37.555 59.115 37.725 69.155 ;
        RECT 39.135 59.115 39.305 69.155 ;
        RECT 40.715 59.115 40.885 69.155 ;
        RECT 42.295 59.115 42.465 69.155 ;
        RECT 45.775 59.115 45.945 69.155 ;
        RECT 47.355 59.115 47.525 69.155 ;
        RECT 48.935 59.115 49.105 69.155 ;
        RECT 50.515 59.115 50.685 69.155 ;
        RECT 52.095 59.115 52.265 69.155 ;
        RECT 55.575 59.115 55.745 69.155 ;
        RECT 57.155 59.115 57.325 69.155 ;
        RECT 58.735 59.115 58.905 69.155 ;
        RECT 60.315 59.115 60.485 69.155 ;
        RECT 61.895 59.115 62.065 69.155 ;
        RECT 65.375 59.115 65.545 69.155 ;
        RECT 66.955 59.115 67.125 69.155 ;
        RECT 68.535 59.115 68.705 69.155 ;
        RECT 70.115 59.115 70.285 69.155 ;
        RECT 71.695 59.115 71.865 69.155 ;
        RECT 26.035 48.035 26.205 58.075 ;
        RECT 27.615 48.035 27.785 58.075 ;
        RECT 29.195 48.035 29.365 58.075 ;
        RECT 30.775 48.035 30.945 58.075 ;
        RECT 32.355 48.035 32.525 58.075 ;
        RECT 35.975 48.035 36.145 58.075 ;
        RECT 37.555 48.035 37.725 58.075 ;
        RECT 39.135 48.035 39.305 58.075 ;
        RECT 40.715 48.035 40.885 58.075 ;
        RECT 42.295 48.035 42.465 58.075 ;
        RECT 45.775 48.035 45.945 58.075 ;
        RECT 47.355 48.035 47.525 58.075 ;
        RECT 48.935 48.035 49.105 58.075 ;
        RECT 50.515 48.035 50.685 58.075 ;
        RECT 52.095 48.035 52.265 58.075 ;
        RECT 55.575 48.035 55.745 58.075 ;
        RECT 57.155 48.035 57.325 58.075 ;
        RECT 58.735 48.035 58.905 58.075 ;
        RECT 60.315 48.035 60.485 58.075 ;
        RECT 61.895 48.035 62.065 58.075 ;
        RECT 65.375 48.035 65.545 58.075 ;
        RECT 66.955 48.035 67.125 58.075 ;
        RECT 68.535 48.035 68.705 58.075 ;
        RECT 70.115 48.035 70.285 58.075 ;
        RECT 71.695 48.035 71.865 58.075 ;
        RECT 26.030 35.005 26.200 45.045 ;
        RECT 27.610 35.005 27.780 45.045 ;
        RECT 29.190 35.005 29.360 45.045 ;
        RECT 30.770 35.005 30.940 45.045 ;
        RECT 32.350 35.005 32.520 45.045 ;
        RECT 35.970 35.005 36.140 45.045 ;
        RECT 37.550 35.005 37.720 45.045 ;
        RECT 39.130 35.005 39.300 45.045 ;
        RECT 40.710 35.005 40.880 45.045 ;
        RECT 42.290 35.005 42.460 45.045 ;
        RECT 45.770 35.005 45.940 45.045 ;
        RECT 47.350 35.005 47.520 45.045 ;
        RECT 48.930 35.005 49.100 45.045 ;
        RECT 50.510 35.005 50.680 45.045 ;
        RECT 52.090 35.005 52.260 45.045 ;
        RECT 55.570 35.005 55.740 45.045 ;
        RECT 57.150 35.005 57.320 45.045 ;
        RECT 58.730 35.005 58.900 45.045 ;
        RECT 60.310 35.005 60.480 45.045 ;
        RECT 61.890 35.005 62.060 45.045 ;
        RECT 65.370 35.005 65.540 45.045 ;
        RECT 66.950 35.005 67.120 45.045 ;
        RECT 68.530 35.005 68.700 45.045 ;
        RECT 70.110 35.005 70.280 45.045 ;
        RECT 71.690 35.005 71.860 45.045 ;
        RECT 26.030 23.825 26.200 33.865 ;
        RECT 27.610 23.825 27.780 33.865 ;
        RECT 29.190 23.825 29.360 33.865 ;
        RECT 30.770 23.825 30.940 33.865 ;
        RECT 32.350 23.825 32.520 33.865 ;
        RECT 35.970 23.825 36.140 33.865 ;
        RECT 37.550 23.825 37.720 33.865 ;
        RECT 39.130 23.825 39.300 33.865 ;
        RECT 40.710 23.825 40.880 33.865 ;
        RECT 42.290 23.825 42.460 33.865 ;
        RECT 45.770 23.825 45.940 33.865 ;
        RECT 47.350 23.825 47.520 33.865 ;
        RECT 48.930 23.825 49.100 33.865 ;
        RECT 50.510 23.825 50.680 33.865 ;
        RECT 52.090 23.825 52.260 33.865 ;
        RECT 55.570 23.825 55.740 33.865 ;
        RECT 57.150 23.825 57.320 33.865 ;
        RECT 58.730 23.825 58.900 33.865 ;
        RECT 60.310 23.825 60.480 33.865 ;
        RECT 61.890 23.825 62.060 33.865 ;
        RECT 65.370 23.825 65.540 33.865 ;
        RECT 66.950 23.825 67.120 33.865 ;
        RECT 68.530 23.825 68.700 33.865 ;
        RECT 70.110 23.825 70.280 33.865 ;
        RECT 71.690 23.825 71.860 33.865 ;
        RECT 26.030 12.645 26.200 22.685 ;
        RECT 27.610 12.645 27.780 22.685 ;
        RECT 29.190 12.645 29.360 22.685 ;
        RECT 30.770 12.645 30.940 22.685 ;
        RECT 32.350 12.645 32.520 22.685 ;
        RECT 35.970 12.645 36.140 22.685 ;
        RECT 37.550 12.645 37.720 22.685 ;
        RECT 39.130 12.645 39.300 22.685 ;
        RECT 40.710 12.645 40.880 22.685 ;
        RECT 42.290 12.645 42.460 22.685 ;
        RECT 45.770 12.645 45.940 22.685 ;
        RECT 47.350 12.645 47.520 22.685 ;
        RECT 48.930 12.645 49.100 22.685 ;
        RECT 50.510 12.645 50.680 22.685 ;
        RECT 52.090 12.645 52.260 22.685 ;
        RECT 55.570 12.645 55.740 22.685 ;
        RECT 57.150 12.645 57.320 22.685 ;
        RECT 58.730 12.645 58.900 22.685 ;
        RECT 60.310 12.645 60.480 22.685 ;
        RECT 61.890 12.645 62.060 22.685 ;
        RECT 65.370 12.645 65.540 22.685 ;
        RECT 66.950 12.645 67.120 22.685 ;
        RECT 68.530 12.645 68.700 22.685 ;
        RECT 70.110 12.645 70.280 22.685 ;
        RECT 71.690 12.645 71.860 22.685 ;
        RECT 26.030 1.465 26.200 11.505 ;
        RECT 27.610 1.465 27.780 11.505 ;
        RECT 29.190 1.465 29.360 11.505 ;
        RECT 30.770 1.465 30.940 11.505 ;
        RECT 32.350 1.465 32.520 11.505 ;
        RECT 35.970 1.465 36.140 11.505 ;
        RECT 37.550 1.465 37.720 11.505 ;
        RECT 39.130 1.465 39.300 11.505 ;
        RECT 40.710 1.465 40.880 11.505 ;
        RECT 42.290 1.465 42.460 11.505 ;
        RECT 45.770 1.465 45.940 11.505 ;
        RECT 47.350 1.465 47.520 11.505 ;
        RECT 48.930 1.465 49.100 11.505 ;
        RECT 50.510 1.465 50.680 11.505 ;
        RECT 52.090 1.465 52.260 11.505 ;
        RECT 55.570 1.465 55.740 11.505 ;
        RECT 57.150 1.465 57.320 11.505 ;
        RECT 58.730 1.465 58.900 11.505 ;
        RECT 60.310 1.465 60.480 11.505 ;
        RECT 61.890 1.465 62.060 11.505 ;
        RECT 65.370 1.465 65.540 11.505 ;
        RECT 66.950 1.465 67.120 11.505 ;
        RECT 68.530 1.465 68.700 11.505 ;
        RECT 70.110 1.465 70.280 11.505 ;
        RECT 71.690 1.465 71.860 11.505 ;
      LAYER mcon ;
        RECT 26.035 59.195 26.205 69.075 ;
        RECT 27.615 59.195 27.785 69.075 ;
        RECT 29.195 59.195 29.365 69.075 ;
        RECT 30.775 59.195 30.945 69.075 ;
        RECT 32.355 59.195 32.525 69.075 ;
        RECT 35.975 59.195 36.145 69.075 ;
        RECT 37.555 59.195 37.725 69.075 ;
        RECT 39.135 59.195 39.305 69.075 ;
        RECT 40.715 59.195 40.885 69.075 ;
        RECT 42.295 59.195 42.465 69.075 ;
        RECT 45.775 59.195 45.945 69.075 ;
        RECT 47.355 59.195 47.525 69.075 ;
        RECT 48.935 59.195 49.105 69.075 ;
        RECT 50.515 59.195 50.685 69.075 ;
        RECT 52.095 59.195 52.265 69.075 ;
        RECT 55.575 59.195 55.745 69.075 ;
        RECT 57.155 59.195 57.325 69.075 ;
        RECT 58.735 59.195 58.905 69.075 ;
        RECT 60.315 59.195 60.485 69.075 ;
        RECT 61.895 59.195 62.065 69.075 ;
        RECT 65.375 59.195 65.545 69.075 ;
        RECT 66.955 59.195 67.125 69.075 ;
        RECT 68.535 59.195 68.705 69.075 ;
        RECT 70.115 59.195 70.285 69.075 ;
        RECT 71.695 59.195 71.865 69.075 ;
        RECT 26.035 48.115 26.205 57.995 ;
        RECT 27.615 48.115 27.785 57.995 ;
        RECT 29.195 48.115 29.365 57.995 ;
        RECT 30.775 48.115 30.945 57.995 ;
        RECT 32.355 48.115 32.525 57.995 ;
        RECT 35.975 48.115 36.145 57.995 ;
        RECT 37.555 48.115 37.725 57.995 ;
        RECT 39.135 48.115 39.305 57.995 ;
        RECT 40.715 48.115 40.885 57.995 ;
        RECT 42.295 48.115 42.465 57.995 ;
        RECT 45.775 48.115 45.945 57.995 ;
        RECT 47.355 48.115 47.525 57.995 ;
        RECT 48.935 48.115 49.105 57.995 ;
        RECT 50.515 48.115 50.685 57.995 ;
        RECT 52.095 48.115 52.265 57.995 ;
        RECT 55.575 48.115 55.745 57.995 ;
        RECT 57.155 48.115 57.325 57.995 ;
        RECT 58.735 48.115 58.905 57.995 ;
        RECT 60.315 48.115 60.485 57.995 ;
        RECT 61.895 48.115 62.065 57.995 ;
        RECT 65.375 48.115 65.545 57.995 ;
        RECT 66.955 48.115 67.125 57.995 ;
        RECT 68.535 48.115 68.705 57.995 ;
        RECT 70.115 48.115 70.285 57.995 ;
        RECT 71.695 48.115 71.865 57.995 ;
        RECT 26.030 35.085 26.200 44.965 ;
        RECT 27.610 35.085 27.780 44.965 ;
        RECT 29.190 35.085 29.360 44.965 ;
        RECT 30.770 35.085 30.940 44.965 ;
        RECT 32.350 35.085 32.520 44.965 ;
        RECT 35.970 35.085 36.140 44.965 ;
        RECT 37.550 35.085 37.720 44.965 ;
        RECT 39.130 35.085 39.300 44.965 ;
        RECT 40.710 35.085 40.880 44.965 ;
        RECT 42.290 35.085 42.460 44.965 ;
        RECT 45.770 35.085 45.940 44.965 ;
        RECT 47.350 35.085 47.520 44.965 ;
        RECT 48.930 35.085 49.100 44.965 ;
        RECT 50.510 35.085 50.680 44.965 ;
        RECT 52.090 35.085 52.260 44.965 ;
        RECT 55.570 35.085 55.740 44.965 ;
        RECT 57.150 35.085 57.320 44.965 ;
        RECT 58.730 35.085 58.900 44.965 ;
        RECT 60.310 35.085 60.480 44.965 ;
        RECT 61.890 35.085 62.060 44.965 ;
        RECT 65.370 35.085 65.540 44.965 ;
        RECT 66.950 35.085 67.120 44.965 ;
        RECT 68.530 35.085 68.700 44.965 ;
        RECT 70.110 35.085 70.280 44.965 ;
        RECT 71.690 35.085 71.860 44.965 ;
        RECT 26.030 23.905 26.200 33.785 ;
        RECT 27.610 23.905 27.780 33.785 ;
        RECT 29.190 23.905 29.360 33.785 ;
        RECT 30.770 23.905 30.940 33.785 ;
        RECT 32.350 23.905 32.520 33.785 ;
        RECT 35.970 23.905 36.140 33.785 ;
        RECT 37.550 23.905 37.720 33.785 ;
        RECT 39.130 23.905 39.300 33.785 ;
        RECT 40.710 23.905 40.880 33.785 ;
        RECT 42.290 23.905 42.460 33.785 ;
        RECT 45.770 23.905 45.940 33.785 ;
        RECT 47.350 23.905 47.520 33.785 ;
        RECT 48.930 23.905 49.100 33.785 ;
        RECT 50.510 23.905 50.680 33.785 ;
        RECT 52.090 23.905 52.260 33.785 ;
        RECT 55.570 23.905 55.740 33.785 ;
        RECT 57.150 23.905 57.320 33.785 ;
        RECT 58.730 23.905 58.900 33.785 ;
        RECT 60.310 23.905 60.480 33.785 ;
        RECT 61.890 23.905 62.060 33.785 ;
        RECT 65.370 23.905 65.540 33.785 ;
        RECT 66.950 23.905 67.120 33.785 ;
        RECT 68.530 23.905 68.700 33.785 ;
        RECT 70.110 23.905 70.280 33.785 ;
        RECT 71.690 23.905 71.860 33.785 ;
        RECT 26.030 12.725 26.200 22.605 ;
        RECT 27.610 12.725 27.780 22.605 ;
        RECT 29.190 12.725 29.360 22.605 ;
        RECT 30.770 12.725 30.940 22.605 ;
        RECT 32.350 12.725 32.520 22.605 ;
        RECT 35.970 12.725 36.140 22.605 ;
        RECT 37.550 12.725 37.720 22.605 ;
        RECT 39.130 12.725 39.300 22.605 ;
        RECT 40.710 12.725 40.880 22.605 ;
        RECT 42.290 12.725 42.460 22.605 ;
        RECT 45.770 12.725 45.940 22.605 ;
        RECT 47.350 12.725 47.520 22.605 ;
        RECT 48.930 12.725 49.100 22.605 ;
        RECT 50.510 12.725 50.680 22.605 ;
        RECT 52.090 12.725 52.260 22.605 ;
        RECT 55.570 12.725 55.740 22.605 ;
        RECT 57.150 12.725 57.320 22.605 ;
        RECT 58.730 12.725 58.900 22.605 ;
        RECT 60.310 12.725 60.480 22.605 ;
        RECT 61.890 12.725 62.060 22.605 ;
        RECT 65.370 12.725 65.540 22.605 ;
        RECT 66.950 12.725 67.120 22.605 ;
        RECT 68.530 12.725 68.700 22.605 ;
        RECT 70.110 12.725 70.280 22.605 ;
        RECT 71.690 12.725 71.860 22.605 ;
        RECT 26.030 1.545 26.200 11.425 ;
        RECT 27.610 1.545 27.780 11.425 ;
        RECT 29.190 1.545 29.360 11.425 ;
        RECT 30.770 1.545 30.940 11.425 ;
        RECT 32.350 1.545 32.520 11.425 ;
        RECT 35.970 1.545 36.140 11.425 ;
        RECT 37.550 1.545 37.720 11.425 ;
        RECT 39.130 1.545 39.300 11.425 ;
        RECT 40.710 1.545 40.880 11.425 ;
        RECT 42.290 1.545 42.460 11.425 ;
        RECT 45.770 1.545 45.940 11.425 ;
        RECT 47.350 1.545 47.520 11.425 ;
        RECT 48.930 1.545 49.100 11.425 ;
        RECT 50.510 1.545 50.680 11.425 ;
        RECT 52.090 1.545 52.260 11.425 ;
        RECT 55.570 1.545 55.740 11.425 ;
        RECT 57.150 1.545 57.320 11.425 ;
        RECT 58.730 1.545 58.900 11.425 ;
        RECT 60.310 1.545 60.480 11.425 ;
        RECT 61.890 1.545 62.060 11.425 ;
        RECT 65.370 1.545 65.540 11.425 ;
        RECT 66.950 1.545 67.120 11.425 ;
        RECT 68.530 1.545 68.700 11.425 ;
        RECT 70.110 1.545 70.280 11.425 ;
        RECT 71.690 1.545 71.860 11.425 ;
      LAYER met1 ;
        RECT 26.005 63.920 26.235 69.135 ;
        RECT 27.585 63.920 27.815 69.135 ;
        RECT 29.165 63.930 29.395 69.135 ;
        RECT 30.745 63.930 30.975 69.135 ;
        RECT 32.325 63.930 32.555 69.135 ;
        RECT 25.730 59.570 26.460 63.920 ;
        RECT 27.320 59.570 28.050 63.920 ;
        RECT 28.890 59.580 29.620 63.930 ;
        RECT 30.470 59.580 31.200 63.930 ;
        RECT 32.060 59.580 32.790 63.930 ;
        RECT 35.945 63.920 36.175 69.135 ;
        RECT 37.525 63.920 37.755 69.135 ;
        RECT 39.105 63.930 39.335 69.135 ;
        RECT 40.685 63.930 40.915 69.135 ;
        RECT 42.265 63.930 42.495 69.135 ;
        RECT 26.005 59.135 26.235 59.570 ;
        RECT 27.585 59.135 27.815 59.570 ;
        RECT 29.165 59.135 29.395 59.580 ;
        RECT 30.745 59.135 30.975 59.580 ;
        RECT 32.325 59.135 32.555 59.580 ;
        RECT 35.660 59.570 36.390 63.920 ;
        RECT 37.250 59.570 37.980 63.920 ;
        RECT 38.820 59.580 39.550 63.930 ;
        RECT 40.400 59.580 41.130 63.930 ;
        RECT 41.990 59.580 42.720 63.930 ;
        RECT 45.745 63.920 45.975 69.135 ;
        RECT 47.325 63.920 47.555 69.135 ;
        RECT 48.905 63.930 49.135 69.135 ;
        RECT 50.485 63.930 50.715 69.135 ;
        RECT 52.065 63.930 52.295 69.135 ;
        RECT 55.545 63.950 55.775 69.135 ;
        RECT 57.125 63.950 57.355 69.135 ;
        RECT 58.705 63.960 58.935 69.135 ;
        RECT 60.285 63.960 60.515 69.135 ;
        RECT 61.865 63.960 62.095 69.135 ;
        RECT 35.945 59.135 36.175 59.570 ;
        RECT 37.525 59.135 37.755 59.570 ;
        RECT 39.105 59.135 39.335 59.580 ;
        RECT 40.685 59.135 40.915 59.580 ;
        RECT 42.265 59.135 42.495 59.580 ;
        RECT 45.470 59.570 46.200 63.920 ;
        RECT 47.060 59.570 47.790 63.920 ;
        RECT 48.630 59.580 49.360 63.930 ;
        RECT 50.210 59.580 50.940 63.930 ;
        RECT 51.800 59.580 52.530 63.930 ;
        RECT 55.280 59.600 56.010 63.950 ;
        RECT 56.870 59.600 57.600 63.950 ;
        RECT 58.440 59.610 59.170 63.960 ;
        RECT 60.020 59.610 60.750 63.960 ;
        RECT 61.610 59.610 62.340 63.960 ;
        RECT 65.345 63.950 65.575 69.135 ;
        RECT 66.925 63.950 67.155 69.135 ;
        RECT 68.505 63.960 68.735 69.135 ;
        RECT 70.085 63.960 70.315 69.135 ;
        RECT 71.665 63.960 71.895 69.135 ;
        RECT 45.745 59.135 45.975 59.570 ;
        RECT 47.325 59.135 47.555 59.570 ;
        RECT 48.905 59.135 49.135 59.580 ;
        RECT 50.485 59.135 50.715 59.580 ;
        RECT 52.065 59.135 52.295 59.580 ;
        RECT 55.545 59.135 55.775 59.600 ;
        RECT 57.125 59.135 57.355 59.600 ;
        RECT 58.705 59.135 58.935 59.610 ;
        RECT 60.285 59.135 60.515 59.610 ;
        RECT 61.865 59.135 62.095 59.610 ;
        RECT 65.070 59.600 65.800 63.950 ;
        RECT 66.660 59.600 67.390 63.950 ;
        RECT 68.230 59.610 68.960 63.960 ;
        RECT 69.810 59.610 70.540 63.960 ;
        RECT 71.400 59.610 72.130 63.960 ;
        RECT 65.345 59.135 65.575 59.600 ;
        RECT 66.925 59.135 67.155 59.600 ;
        RECT 68.505 59.135 68.735 59.610 ;
        RECT 70.085 59.135 70.315 59.610 ;
        RECT 71.665 59.135 71.895 59.610 ;
        RECT 26.005 52.870 26.235 58.055 ;
        RECT 27.585 52.870 27.815 58.055 ;
        RECT 29.165 52.880 29.395 58.055 ;
        RECT 30.745 52.880 30.975 58.055 ;
        RECT 32.325 52.880 32.555 58.055 ;
        RECT 25.720 48.520 26.450 52.870 ;
        RECT 27.310 48.520 28.040 52.870 ;
        RECT 28.880 48.530 29.610 52.880 ;
        RECT 30.460 48.530 31.190 52.880 ;
        RECT 32.050 48.530 32.780 52.880 ;
        RECT 35.945 52.870 36.175 58.055 ;
        RECT 37.525 52.870 37.755 58.055 ;
        RECT 39.105 52.880 39.335 58.055 ;
        RECT 40.685 52.880 40.915 58.055 ;
        RECT 42.265 52.880 42.495 58.055 ;
        RECT 26.005 48.055 26.235 48.520 ;
        RECT 27.585 48.055 27.815 48.520 ;
        RECT 29.165 48.055 29.395 48.530 ;
        RECT 30.745 48.055 30.975 48.530 ;
        RECT 32.325 48.055 32.555 48.530 ;
        RECT 35.650 48.520 36.380 52.870 ;
        RECT 37.240 48.520 37.970 52.870 ;
        RECT 38.810 48.530 39.540 52.880 ;
        RECT 40.390 48.530 41.120 52.880 ;
        RECT 41.980 48.530 42.710 52.880 ;
        RECT 45.745 52.870 45.975 58.055 ;
        RECT 47.325 52.870 47.555 58.055 ;
        RECT 48.905 52.880 49.135 58.055 ;
        RECT 50.485 52.880 50.715 58.055 ;
        RECT 52.065 52.880 52.295 58.055 ;
        RECT 55.545 52.900 55.775 58.055 ;
        RECT 57.125 52.900 57.355 58.055 ;
        RECT 58.705 52.910 58.935 58.055 ;
        RECT 60.285 52.910 60.515 58.055 ;
        RECT 61.865 52.910 62.095 58.055 ;
        RECT 35.945 48.055 36.175 48.520 ;
        RECT 37.525 48.055 37.755 48.520 ;
        RECT 39.105 48.055 39.335 48.530 ;
        RECT 40.685 48.055 40.915 48.530 ;
        RECT 42.265 48.055 42.495 48.530 ;
        RECT 45.460 48.520 46.190 52.870 ;
        RECT 47.050 48.520 47.780 52.870 ;
        RECT 48.620 48.530 49.350 52.880 ;
        RECT 50.200 48.530 50.930 52.880 ;
        RECT 51.790 48.530 52.520 52.880 ;
        RECT 55.270 48.550 56.000 52.900 ;
        RECT 56.860 48.550 57.590 52.900 ;
        RECT 58.430 48.560 59.160 52.910 ;
        RECT 60.010 48.560 60.740 52.910 ;
        RECT 61.600 48.560 62.330 52.910 ;
        RECT 65.345 52.900 65.575 58.055 ;
        RECT 66.925 52.900 67.155 58.055 ;
        RECT 68.505 52.910 68.735 58.055 ;
        RECT 70.085 52.910 70.315 58.055 ;
        RECT 71.665 52.910 71.895 58.055 ;
        RECT 45.745 48.055 45.975 48.520 ;
        RECT 47.325 48.055 47.555 48.520 ;
        RECT 48.905 48.055 49.135 48.530 ;
        RECT 50.485 48.055 50.715 48.530 ;
        RECT 52.065 48.055 52.295 48.530 ;
        RECT 55.545 48.055 55.775 48.550 ;
        RECT 57.125 48.055 57.355 48.550 ;
        RECT 58.705 48.055 58.935 48.560 ;
        RECT 60.285 48.055 60.515 48.560 ;
        RECT 61.865 48.055 62.095 48.560 ;
        RECT 65.060 48.550 65.790 52.900 ;
        RECT 66.650 48.550 67.380 52.900 ;
        RECT 68.220 48.560 68.950 52.910 ;
        RECT 69.800 48.560 70.530 52.910 ;
        RECT 71.390 48.560 72.120 52.910 ;
        RECT 65.345 48.055 65.575 48.550 ;
        RECT 66.925 48.055 67.155 48.550 ;
        RECT 68.505 48.055 68.735 48.560 ;
        RECT 70.085 48.055 70.315 48.560 ;
        RECT 71.665 48.055 71.895 48.560 ;
        RECT 26.000 39.840 26.230 45.025 ;
        RECT 27.580 39.840 27.810 45.025 ;
        RECT 29.160 39.850 29.390 45.025 ;
        RECT 30.740 39.850 30.970 45.025 ;
        RECT 32.320 39.850 32.550 45.025 ;
        RECT 25.720 35.490 26.450 39.840 ;
        RECT 27.310 35.490 28.040 39.840 ;
        RECT 28.880 35.500 29.610 39.850 ;
        RECT 30.460 35.500 31.190 39.850 ;
        RECT 32.050 35.500 32.780 39.850 ;
        RECT 35.940 39.840 36.170 45.025 ;
        RECT 37.520 39.840 37.750 45.025 ;
        RECT 39.100 39.850 39.330 45.025 ;
        RECT 40.680 39.850 40.910 45.025 ;
        RECT 42.260 39.850 42.490 45.025 ;
        RECT 26.000 35.025 26.230 35.490 ;
        RECT 27.580 35.025 27.810 35.490 ;
        RECT 29.160 35.025 29.390 35.500 ;
        RECT 30.740 35.025 30.970 35.500 ;
        RECT 32.320 35.025 32.550 35.500 ;
        RECT 35.650 35.490 36.380 39.840 ;
        RECT 37.240 35.490 37.970 39.840 ;
        RECT 38.810 35.500 39.540 39.850 ;
        RECT 40.390 35.500 41.120 39.850 ;
        RECT 41.980 35.500 42.710 39.850 ;
        RECT 45.740 39.840 45.970 45.025 ;
        RECT 47.320 39.840 47.550 45.025 ;
        RECT 48.900 39.850 49.130 45.025 ;
        RECT 50.480 39.850 50.710 45.025 ;
        RECT 52.060 39.850 52.290 45.025 ;
        RECT 55.540 39.870 55.770 45.025 ;
        RECT 57.120 39.870 57.350 45.025 ;
        RECT 58.700 39.880 58.930 45.025 ;
        RECT 60.280 39.880 60.510 45.025 ;
        RECT 61.860 39.880 62.090 45.025 ;
        RECT 35.940 35.025 36.170 35.490 ;
        RECT 37.520 35.025 37.750 35.490 ;
        RECT 39.100 35.025 39.330 35.500 ;
        RECT 40.680 35.025 40.910 35.500 ;
        RECT 42.260 35.025 42.490 35.500 ;
        RECT 45.460 35.490 46.190 39.840 ;
        RECT 47.050 35.490 47.780 39.840 ;
        RECT 48.620 35.500 49.350 39.850 ;
        RECT 50.200 35.500 50.930 39.850 ;
        RECT 51.790 35.500 52.520 39.850 ;
        RECT 55.270 35.520 56.000 39.870 ;
        RECT 56.860 35.520 57.590 39.870 ;
        RECT 58.430 35.530 59.160 39.880 ;
        RECT 60.010 35.530 60.740 39.880 ;
        RECT 61.600 35.530 62.330 39.880 ;
        RECT 65.340 39.870 65.570 45.025 ;
        RECT 66.920 39.870 67.150 45.025 ;
        RECT 68.500 39.880 68.730 45.025 ;
        RECT 70.080 39.880 70.310 45.025 ;
        RECT 71.660 39.880 71.890 45.025 ;
        RECT 45.740 35.025 45.970 35.490 ;
        RECT 47.320 35.025 47.550 35.490 ;
        RECT 48.900 35.025 49.130 35.500 ;
        RECT 50.480 35.025 50.710 35.500 ;
        RECT 52.060 35.025 52.290 35.500 ;
        RECT 55.540 35.025 55.770 35.520 ;
        RECT 57.120 35.025 57.350 35.520 ;
        RECT 58.700 35.025 58.930 35.530 ;
        RECT 60.280 35.025 60.510 35.530 ;
        RECT 61.860 35.025 62.090 35.530 ;
        RECT 65.060 35.520 65.790 39.870 ;
        RECT 66.650 35.520 67.380 39.870 ;
        RECT 68.220 35.530 68.950 39.880 ;
        RECT 69.800 35.530 70.530 39.880 ;
        RECT 71.390 35.530 72.120 39.880 ;
        RECT 65.340 35.025 65.570 35.520 ;
        RECT 66.920 35.025 67.150 35.520 ;
        RECT 68.500 35.025 68.730 35.530 ;
        RECT 70.080 35.025 70.310 35.530 ;
        RECT 71.660 35.025 71.890 35.530 ;
        RECT 26.000 28.660 26.230 33.845 ;
        RECT 27.580 28.660 27.810 33.845 ;
        RECT 29.160 28.670 29.390 33.845 ;
        RECT 30.740 28.670 30.970 33.845 ;
        RECT 32.320 28.670 32.550 33.845 ;
        RECT 25.720 24.310 26.450 28.660 ;
        RECT 27.310 24.310 28.040 28.660 ;
        RECT 28.880 24.320 29.610 28.670 ;
        RECT 30.460 24.320 31.190 28.670 ;
        RECT 32.050 24.320 32.780 28.670 ;
        RECT 35.940 28.660 36.170 33.845 ;
        RECT 37.520 28.660 37.750 33.845 ;
        RECT 39.100 28.670 39.330 33.845 ;
        RECT 40.680 28.670 40.910 33.845 ;
        RECT 42.260 28.670 42.490 33.845 ;
        RECT 26.000 23.845 26.230 24.310 ;
        RECT 27.580 23.845 27.810 24.310 ;
        RECT 29.160 23.845 29.390 24.320 ;
        RECT 30.740 23.845 30.970 24.320 ;
        RECT 32.320 23.845 32.550 24.320 ;
        RECT 35.650 24.310 36.380 28.660 ;
        RECT 37.240 24.310 37.970 28.660 ;
        RECT 38.810 24.320 39.540 28.670 ;
        RECT 40.390 24.320 41.120 28.670 ;
        RECT 41.980 24.320 42.710 28.670 ;
        RECT 45.740 28.660 45.970 33.845 ;
        RECT 47.320 28.660 47.550 33.845 ;
        RECT 48.900 28.670 49.130 33.845 ;
        RECT 50.480 28.670 50.710 33.845 ;
        RECT 52.060 28.670 52.290 33.845 ;
        RECT 55.540 28.690 55.770 33.845 ;
        RECT 57.120 28.690 57.350 33.845 ;
        RECT 58.700 28.700 58.930 33.845 ;
        RECT 60.280 28.700 60.510 33.845 ;
        RECT 61.860 28.700 62.090 33.845 ;
        RECT 35.940 23.845 36.170 24.310 ;
        RECT 37.520 23.845 37.750 24.310 ;
        RECT 39.100 23.845 39.330 24.320 ;
        RECT 40.680 23.845 40.910 24.320 ;
        RECT 42.260 23.845 42.490 24.320 ;
        RECT 45.460 24.310 46.190 28.660 ;
        RECT 47.050 24.310 47.780 28.660 ;
        RECT 48.620 24.320 49.350 28.670 ;
        RECT 50.200 24.320 50.930 28.670 ;
        RECT 51.790 24.320 52.520 28.670 ;
        RECT 55.270 24.340 56.000 28.690 ;
        RECT 56.860 24.340 57.590 28.690 ;
        RECT 58.430 24.350 59.160 28.700 ;
        RECT 60.010 24.350 60.740 28.700 ;
        RECT 61.600 24.350 62.330 28.700 ;
        RECT 65.340 28.690 65.570 33.845 ;
        RECT 66.920 28.690 67.150 33.845 ;
        RECT 68.500 28.700 68.730 33.845 ;
        RECT 70.080 28.700 70.310 33.845 ;
        RECT 71.660 28.700 71.890 33.845 ;
        RECT 45.740 23.845 45.970 24.310 ;
        RECT 47.320 23.845 47.550 24.310 ;
        RECT 48.900 23.845 49.130 24.320 ;
        RECT 50.480 23.845 50.710 24.320 ;
        RECT 52.060 23.845 52.290 24.320 ;
        RECT 55.540 23.845 55.770 24.340 ;
        RECT 57.120 23.845 57.350 24.340 ;
        RECT 58.700 23.845 58.930 24.350 ;
        RECT 60.280 23.845 60.510 24.350 ;
        RECT 61.860 23.845 62.090 24.350 ;
        RECT 65.060 24.340 65.790 28.690 ;
        RECT 66.650 24.340 67.380 28.690 ;
        RECT 68.220 24.350 68.950 28.700 ;
        RECT 69.800 24.350 70.530 28.700 ;
        RECT 71.390 24.350 72.120 28.700 ;
        RECT 65.340 23.845 65.570 24.340 ;
        RECT 66.920 23.845 67.150 24.340 ;
        RECT 68.500 23.845 68.730 24.350 ;
        RECT 70.080 23.845 70.310 24.350 ;
        RECT 71.660 23.845 71.890 24.350 ;
        RECT 26.000 17.480 26.230 22.665 ;
        RECT 27.580 17.480 27.810 22.665 ;
        RECT 29.160 17.490 29.390 22.665 ;
        RECT 30.740 17.490 30.970 22.665 ;
        RECT 32.320 17.490 32.550 22.665 ;
        RECT 25.720 13.130 26.450 17.480 ;
        RECT 27.310 13.130 28.040 17.480 ;
        RECT 28.880 13.140 29.610 17.490 ;
        RECT 30.460 13.140 31.190 17.490 ;
        RECT 32.050 13.140 32.780 17.490 ;
        RECT 35.940 17.480 36.170 22.665 ;
        RECT 37.520 17.480 37.750 22.665 ;
        RECT 39.100 17.490 39.330 22.665 ;
        RECT 40.680 17.490 40.910 22.665 ;
        RECT 42.260 17.490 42.490 22.665 ;
        RECT 26.000 12.665 26.230 13.130 ;
        RECT 27.580 12.665 27.810 13.130 ;
        RECT 29.160 12.665 29.390 13.140 ;
        RECT 30.740 12.665 30.970 13.140 ;
        RECT 32.320 12.665 32.550 13.140 ;
        RECT 35.650 13.130 36.380 17.480 ;
        RECT 37.240 13.130 37.970 17.480 ;
        RECT 38.810 13.140 39.540 17.490 ;
        RECT 40.390 13.140 41.120 17.490 ;
        RECT 41.980 13.140 42.710 17.490 ;
        RECT 45.740 17.480 45.970 22.665 ;
        RECT 47.320 17.480 47.550 22.665 ;
        RECT 48.900 17.490 49.130 22.665 ;
        RECT 50.480 17.490 50.710 22.665 ;
        RECT 52.060 17.490 52.290 22.665 ;
        RECT 55.540 17.510 55.770 22.665 ;
        RECT 57.120 17.510 57.350 22.665 ;
        RECT 58.700 17.520 58.930 22.665 ;
        RECT 60.280 17.520 60.510 22.665 ;
        RECT 61.860 17.520 62.090 22.665 ;
        RECT 35.940 12.665 36.170 13.130 ;
        RECT 37.520 12.665 37.750 13.130 ;
        RECT 39.100 12.665 39.330 13.140 ;
        RECT 40.680 12.665 40.910 13.140 ;
        RECT 42.260 12.665 42.490 13.140 ;
        RECT 45.460 13.130 46.190 17.480 ;
        RECT 47.050 13.130 47.780 17.480 ;
        RECT 48.620 13.140 49.350 17.490 ;
        RECT 50.200 13.140 50.930 17.490 ;
        RECT 51.790 13.140 52.520 17.490 ;
        RECT 55.270 13.160 56.000 17.510 ;
        RECT 56.860 13.160 57.590 17.510 ;
        RECT 58.430 13.170 59.160 17.520 ;
        RECT 60.010 13.170 60.740 17.520 ;
        RECT 61.600 13.170 62.330 17.520 ;
        RECT 65.340 17.510 65.570 22.665 ;
        RECT 66.920 17.510 67.150 22.665 ;
        RECT 68.500 17.520 68.730 22.665 ;
        RECT 70.080 17.520 70.310 22.665 ;
        RECT 71.660 17.520 71.890 22.665 ;
        RECT 45.740 12.665 45.970 13.130 ;
        RECT 47.320 12.665 47.550 13.130 ;
        RECT 48.900 12.665 49.130 13.140 ;
        RECT 50.480 12.665 50.710 13.140 ;
        RECT 52.060 12.665 52.290 13.140 ;
        RECT 55.540 12.665 55.770 13.160 ;
        RECT 57.120 12.665 57.350 13.160 ;
        RECT 58.700 12.665 58.930 13.170 ;
        RECT 60.280 12.665 60.510 13.170 ;
        RECT 61.860 12.665 62.090 13.170 ;
        RECT 65.060 13.160 65.790 17.510 ;
        RECT 66.650 13.160 67.380 17.510 ;
        RECT 68.220 13.170 68.950 17.520 ;
        RECT 69.800 13.170 70.530 17.520 ;
        RECT 71.390 13.170 72.120 17.520 ;
        RECT 65.340 12.665 65.570 13.160 ;
        RECT 66.920 12.665 67.150 13.160 ;
        RECT 68.500 12.665 68.730 13.170 ;
        RECT 70.080 12.665 70.310 13.170 ;
        RECT 71.660 12.665 71.890 13.170 ;
        RECT 26.000 6.300 26.230 11.485 ;
        RECT 27.580 6.300 27.810 11.485 ;
        RECT 29.160 6.310 29.390 11.485 ;
        RECT 30.740 6.310 30.970 11.485 ;
        RECT 32.320 6.310 32.550 11.485 ;
        RECT 25.720 1.950 26.450 6.300 ;
        RECT 27.310 1.950 28.040 6.300 ;
        RECT 28.880 1.960 29.610 6.310 ;
        RECT 30.460 1.960 31.190 6.310 ;
        RECT 32.050 1.960 32.780 6.310 ;
        RECT 35.940 6.300 36.170 11.485 ;
        RECT 37.520 6.300 37.750 11.485 ;
        RECT 39.100 6.310 39.330 11.485 ;
        RECT 40.680 6.310 40.910 11.485 ;
        RECT 42.260 6.310 42.490 11.485 ;
        RECT 26.000 1.485 26.230 1.950 ;
        RECT 27.580 1.485 27.810 1.950 ;
        RECT 29.160 1.485 29.390 1.960 ;
        RECT 30.740 1.485 30.970 1.960 ;
        RECT 32.320 1.485 32.550 1.960 ;
        RECT 35.650 1.950 36.380 6.300 ;
        RECT 37.240 1.950 37.970 6.300 ;
        RECT 38.810 1.960 39.540 6.310 ;
        RECT 40.390 1.960 41.120 6.310 ;
        RECT 41.980 1.960 42.710 6.310 ;
        RECT 45.740 6.300 45.970 11.485 ;
        RECT 47.320 6.300 47.550 11.485 ;
        RECT 48.900 6.310 49.130 11.485 ;
        RECT 50.480 6.310 50.710 11.485 ;
        RECT 52.060 6.310 52.290 11.485 ;
        RECT 55.540 6.330 55.770 11.485 ;
        RECT 57.120 6.330 57.350 11.485 ;
        RECT 58.700 6.340 58.930 11.485 ;
        RECT 60.280 6.340 60.510 11.485 ;
        RECT 61.860 6.340 62.090 11.485 ;
        RECT 35.940 1.485 36.170 1.950 ;
        RECT 37.520 1.485 37.750 1.950 ;
        RECT 39.100 1.485 39.330 1.960 ;
        RECT 40.680 1.485 40.910 1.960 ;
        RECT 42.260 1.485 42.490 1.960 ;
        RECT 45.460 1.950 46.190 6.300 ;
        RECT 47.050 1.950 47.780 6.300 ;
        RECT 48.620 1.960 49.350 6.310 ;
        RECT 50.200 1.960 50.930 6.310 ;
        RECT 51.790 1.960 52.520 6.310 ;
        RECT 55.270 1.980 56.000 6.330 ;
        RECT 56.860 1.980 57.590 6.330 ;
        RECT 58.430 1.990 59.160 6.340 ;
        RECT 60.010 1.990 60.740 6.340 ;
        RECT 61.600 1.990 62.330 6.340 ;
        RECT 65.340 6.330 65.570 11.485 ;
        RECT 66.920 6.330 67.150 11.485 ;
        RECT 68.500 6.340 68.730 11.485 ;
        RECT 70.080 6.340 70.310 11.485 ;
        RECT 71.660 6.340 71.890 11.485 ;
        RECT 45.740 1.485 45.970 1.950 ;
        RECT 47.320 1.485 47.550 1.950 ;
        RECT 48.900 1.485 49.130 1.960 ;
        RECT 50.480 1.485 50.710 1.960 ;
        RECT 52.060 1.485 52.290 1.960 ;
        RECT 55.540 1.485 55.770 1.980 ;
        RECT 57.120 1.485 57.350 1.980 ;
        RECT 58.700 1.485 58.930 1.990 ;
        RECT 60.280 1.485 60.510 1.990 ;
        RECT 61.860 1.485 62.090 1.990 ;
        RECT 65.060 1.980 65.790 6.330 ;
        RECT 66.650 1.980 67.380 6.330 ;
        RECT 68.220 1.990 68.950 6.340 ;
        RECT 69.800 1.990 70.530 6.340 ;
        RECT 71.390 1.990 72.120 6.340 ;
        RECT 65.340 1.485 65.570 1.980 ;
        RECT 66.920 1.485 67.150 1.980 ;
        RECT 68.500 1.485 68.730 1.990 ;
        RECT 70.080 1.485 70.310 1.990 ;
        RECT 71.660 1.485 71.890 1.990 ;
      LAYER via ;
        RECT 25.780 59.570 26.410 63.920 ;
        RECT 27.370 59.570 28.000 63.920 ;
        RECT 28.940 59.580 29.570 63.930 ;
        RECT 30.520 59.580 31.150 63.930 ;
        RECT 32.110 59.580 32.740 63.930 ;
        RECT 35.710 59.570 36.340 63.920 ;
        RECT 37.300 59.570 37.930 63.920 ;
        RECT 38.870 59.580 39.500 63.930 ;
        RECT 40.450 59.580 41.080 63.930 ;
        RECT 42.040 59.580 42.670 63.930 ;
        RECT 45.520 59.570 46.150 63.920 ;
        RECT 47.110 59.570 47.740 63.920 ;
        RECT 48.680 59.580 49.310 63.930 ;
        RECT 50.260 59.580 50.890 63.930 ;
        RECT 51.850 59.580 52.480 63.930 ;
        RECT 55.330 59.600 55.960 63.950 ;
        RECT 56.920 59.600 57.550 63.950 ;
        RECT 58.490 59.610 59.120 63.960 ;
        RECT 60.070 59.610 60.700 63.960 ;
        RECT 61.660 59.610 62.290 63.960 ;
        RECT 65.120 59.600 65.750 63.950 ;
        RECT 66.710 59.600 67.340 63.950 ;
        RECT 68.280 59.610 68.910 63.960 ;
        RECT 69.860 59.610 70.490 63.960 ;
        RECT 71.450 59.610 72.080 63.960 ;
        RECT 25.770 48.520 26.400 52.870 ;
        RECT 27.360 48.520 27.990 52.870 ;
        RECT 28.930 48.530 29.560 52.880 ;
        RECT 30.510 48.530 31.140 52.880 ;
        RECT 32.100 48.530 32.730 52.880 ;
        RECT 35.700 48.520 36.330 52.870 ;
        RECT 37.290 48.520 37.920 52.870 ;
        RECT 38.860 48.530 39.490 52.880 ;
        RECT 40.440 48.530 41.070 52.880 ;
        RECT 42.030 48.530 42.660 52.880 ;
        RECT 45.510 48.520 46.140 52.870 ;
        RECT 47.100 48.520 47.730 52.870 ;
        RECT 48.670 48.530 49.300 52.880 ;
        RECT 50.250 48.530 50.880 52.880 ;
        RECT 51.840 48.530 52.470 52.880 ;
        RECT 55.320 48.550 55.950 52.900 ;
        RECT 56.910 48.550 57.540 52.900 ;
        RECT 58.480 48.560 59.110 52.910 ;
        RECT 60.060 48.560 60.690 52.910 ;
        RECT 61.650 48.560 62.280 52.910 ;
        RECT 65.110 48.550 65.740 52.900 ;
        RECT 66.700 48.550 67.330 52.900 ;
        RECT 68.270 48.560 68.900 52.910 ;
        RECT 69.850 48.560 70.480 52.910 ;
        RECT 71.440 48.560 72.070 52.910 ;
        RECT 25.770 35.490 26.400 39.840 ;
        RECT 27.360 35.490 27.990 39.840 ;
        RECT 28.930 35.500 29.560 39.850 ;
        RECT 30.510 35.500 31.140 39.850 ;
        RECT 32.100 35.500 32.730 39.850 ;
        RECT 35.700 35.490 36.330 39.840 ;
        RECT 37.290 35.490 37.920 39.840 ;
        RECT 38.860 35.500 39.490 39.850 ;
        RECT 40.440 35.500 41.070 39.850 ;
        RECT 42.030 35.500 42.660 39.850 ;
        RECT 45.510 35.490 46.140 39.840 ;
        RECT 47.100 35.490 47.730 39.840 ;
        RECT 48.670 35.500 49.300 39.850 ;
        RECT 50.250 35.500 50.880 39.850 ;
        RECT 51.840 35.500 52.470 39.850 ;
        RECT 55.320 35.520 55.950 39.870 ;
        RECT 56.910 35.520 57.540 39.870 ;
        RECT 58.480 35.530 59.110 39.880 ;
        RECT 60.060 35.530 60.690 39.880 ;
        RECT 61.650 35.530 62.280 39.880 ;
        RECT 65.110 35.520 65.740 39.870 ;
        RECT 66.700 35.520 67.330 39.870 ;
        RECT 68.270 35.530 68.900 39.880 ;
        RECT 69.850 35.530 70.480 39.880 ;
        RECT 71.440 35.530 72.070 39.880 ;
        RECT 25.770 24.310 26.400 28.660 ;
        RECT 27.360 24.310 27.990 28.660 ;
        RECT 28.930 24.320 29.560 28.670 ;
        RECT 30.510 24.320 31.140 28.670 ;
        RECT 32.100 24.320 32.730 28.670 ;
        RECT 35.700 24.310 36.330 28.660 ;
        RECT 37.290 24.310 37.920 28.660 ;
        RECT 38.860 24.320 39.490 28.670 ;
        RECT 40.440 24.320 41.070 28.670 ;
        RECT 42.030 24.320 42.660 28.670 ;
        RECT 45.510 24.310 46.140 28.660 ;
        RECT 47.100 24.310 47.730 28.660 ;
        RECT 48.670 24.320 49.300 28.670 ;
        RECT 50.250 24.320 50.880 28.670 ;
        RECT 51.840 24.320 52.470 28.670 ;
        RECT 55.320 24.340 55.950 28.690 ;
        RECT 56.910 24.340 57.540 28.690 ;
        RECT 58.480 24.350 59.110 28.700 ;
        RECT 60.060 24.350 60.690 28.700 ;
        RECT 61.650 24.350 62.280 28.700 ;
        RECT 65.110 24.340 65.740 28.690 ;
        RECT 66.700 24.340 67.330 28.690 ;
        RECT 68.270 24.350 68.900 28.700 ;
        RECT 69.850 24.350 70.480 28.700 ;
        RECT 71.440 24.350 72.070 28.700 ;
        RECT 25.770 13.130 26.400 17.480 ;
        RECT 27.360 13.130 27.990 17.480 ;
        RECT 28.930 13.140 29.560 17.490 ;
        RECT 30.510 13.140 31.140 17.490 ;
        RECT 32.100 13.140 32.730 17.490 ;
        RECT 35.700 13.130 36.330 17.480 ;
        RECT 37.290 13.130 37.920 17.480 ;
        RECT 38.860 13.140 39.490 17.490 ;
        RECT 40.440 13.140 41.070 17.490 ;
        RECT 42.030 13.140 42.660 17.490 ;
        RECT 45.510 13.130 46.140 17.480 ;
        RECT 47.100 13.130 47.730 17.480 ;
        RECT 48.670 13.140 49.300 17.490 ;
        RECT 50.250 13.140 50.880 17.490 ;
        RECT 51.840 13.140 52.470 17.490 ;
        RECT 55.320 13.160 55.950 17.510 ;
        RECT 56.910 13.160 57.540 17.510 ;
        RECT 58.480 13.170 59.110 17.520 ;
        RECT 60.060 13.170 60.690 17.520 ;
        RECT 61.650 13.170 62.280 17.520 ;
        RECT 65.110 13.160 65.740 17.510 ;
        RECT 66.700 13.160 67.330 17.510 ;
        RECT 68.270 13.170 68.900 17.520 ;
        RECT 69.850 13.170 70.480 17.520 ;
        RECT 71.440 13.170 72.070 17.520 ;
        RECT 25.770 1.950 26.400 6.300 ;
        RECT 27.360 1.950 27.990 6.300 ;
        RECT 28.930 1.960 29.560 6.310 ;
        RECT 30.510 1.960 31.140 6.310 ;
        RECT 32.100 1.960 32.730 6.310 ;
        RECT 35.700 1.950 36.330 6.300 ;
        RECT 37.290 1.950 37.920 6.300 ;
        RECT 38.860 1.960 39.490 6.310 ;
        RECT 40.440 1.960 41.070 6.310 ;
        RECT 42.030 1.960 42.660 6.310 ;
        RECT 45.510 1.950 46.140 6.300 ;
        RECT 47.100 1.950 47.730 6.300 ;
        RECT 48.670 1.960 49.300 6.310 ;
        RECT 50.250 1.960 50.880 6.310 ;
        RECT 51.840 1.960 52.470 6.310 ;
        RECT 55.320 1.980 55.950 6.330 ;
        RECT 56.910 1.980 57.540 6.330 ;
        RECT 58.480 1.990 59.110 6.340 ;
        RECT 60.060 1.990 60.690 6.340 ;
        RECT 61.650 1.990 62.280 6.340 ;
        RECT 65.110 1.980 65.740 6.330 ;
        RECT 66.700 1.980 67.330 6.330 ;
        RECT 68.270 1.990 68.900 6.340 ;
        RECT 69.850 1.990 70.480 6.340 ;
        RECT 71.440 1.990 72.070 6.340 ;
      LAYER met2 ;
        RECT 25.780 63.210 26.410 63.970 ;
        RECT 27.370 63.210 28.000 63.970 ;
        RECT 28.940 63.210 29.570 63.980 ;
        RECT 30.520 63.210 31.150 63.980 ;
        RECT 32.110 63.210 32.740 63.980 ;
        RECT 35.710 63.210 36.340 63.970 ;
        RECT 37.300 63.210 37.930 63.970 ;
        RECT 38.870 63.210 39.500 63.980 ;
        RECT 40.450 63.210 41.080 63.980 ;
        RECT 42.040 63.210 42.670 63.980 ;
        RECT 45.520 63.210 46.150 63.970 ;
        RECT 47.110 63.210 47.740 63.970 ;
        RECT 48.680 63.210 49.310 63.980 ;
        RECT 50.260 63.210 50.890 63.980 ;
        RECT 51.850 63.210 52.480 63.980 ;
        RECT 55.330 63.210 55.960 64.000 ;
        RECT 56.920 63.210 57.550 64.000 ;
        RECT 58.490 63.210 59.120 64.010 ;
        RECT 60.070 63.210 60.700 64.010 ;
        RECT 61.660 63.210 62.290 64.010 ;
        RECT 65.120 63.220 65.750 64.000 ;
        RECT 66.710 63.220 67.340 64.000 ;
        RECT 68.280 63.220 68.910 64.010 ;
        RECT 69.860 63.220 70.490 64.010 ;
        RECT 71.450 63.220 72.080 64.010 ;
        RECT 62.530 63.210 72.080 63.220 ;
        RECT 25.780 60.540 72.080 63.210 ;
        RECT 25.780 59.520 26.410 60.540 ;
        RECT 27.370 59.520 28.000 60.540 ;
        RECT 28.940 59.530 29.570 60.540 ;
        RECT 30.520 59.530 31.150 60.540 ;
        RECT 32.110 59.530 32.740 60.540 ;
        RECT 35.710 59.520 36.340 60.540 ;
        RECT 37.300 59.520 37.930 60.540 ;
        RECT 38.870 59.530 39.500 60.540 ;
        RECT 40.450 59.530 41.080 60.540 ;
        RECT 42.040 59.530 42.670 60.540 ;
        RECT 45.520 59.520 46.150 60.540 ;
        RECT 47.110 59.520 47.740 60.540 ;
        RECT 48.680 59.530 49.310 60.540 ;
        RECT 50.260 59.530 50.890 60.540 ;
        RECT 51.850 59.530 52.480 60.540 ;
        RECT 55.330 59.550 55.960 60.540 ;
        RECT 56.920 59.550 57.550 60.540 ;
        RECT 58.490 59.560 59.120 60.540 ;
        RECT 60.070 59.560 60.700 60.540 ;
        RECT 61.660 59.560 62.290 60.540 ;
        RECT 65.120 59.550 65.750 60.540 ;
        RECT 66.710 59.550 67.340 60.540 ;
        RECT 68.280 59.560 68.910 60.540 ;
        RECT 69.860 59.560 70.490 60.540 ;
        RECT 71.450 59.560 72.080 60.540 ;
        RECT 25.770 51.960 26.400 52.920 ;
        RECT 27.360 51.960 27.990 52.920 ;
        RECT 28.930 51.960 29.560 52.930 ;
        RECT 30.510 51.960 31.140 52.930 ;
        RECT 32.100 51.960 32.730 52.930 ;
        RECT 35.700 51.960 36.330 52.920 ;
        RECT 37.290 51.960 37.920 52.920 ;
        RECT 38.860 51.960 39.490 52.930 ;
        RECT 40.440 51.960 41.070 52.930 ;
        RECT 42.030 51.960 42.660 52.930 ;
        RECT 45.510 51.960 46.140 52.920 ;
        RECT 47.100 51.960 47.730 52.920 ;
        RECT 48.670 51.960 49.300 52.930 ;
        RECT 50.250 51.960 50.880 52.930 ;
        RECT 51.840 51.960 52.470 52.930 ;
        RECT 55.320 51.960 55.950 52.950 ;
        RECT 56.910 51.960 57.540 52.950 ;
        RECT 58.480 51.960 59.110 52.960 ;
        RECT 60.060 51.960 60.690 52.960 ;
        RECT 61.650 51.960 62.280 52.960 ;
        RECT 65.110 51.960 65.740 52.950 ;
        RECT 66.700 51.960 67.330 52.950 ;
        RECT 68.270 51.960 68.900 52.960 ;
        RECT 69.850 51.960 70.480 52.960 ;
        RECT 71.440 51.960 72.070 52.960 ;
        RECT 25.770 49.290 72.070 51.960 ;
        RECT 25.770 48.470 26.400 49.290 ;
        RECT 27.360 48.470 27.990 49.290 ;
        RECT 28.930 48.480 29.560 49.290 ;
        RECT 30.510 48.480 31.140 49.290 ;
        RECT 32.100 48.480 32.730 49.290 ;
        RECT 35.700 48.470 36.330 49.290 ;
        RECT 37.290 48.470 37.920 49.290 ;
        RECT 38.860 48.480 39.490 49.290 ;
        RECT 40.440 48.480 41.070 49.290 ;
        RECT 42.030 48.480 42.660 49.290 ;
        RECT 45.510 48.470 46.140 49.290 ;
        RECT 47.100 48.470 47.730 49.290 ;
        RECT 48.670 48.480 49.300 49.290 ;
        RECT 50.250 48.480 50.880 49.290 ;
        RECT 51.840 48.480 52.470 49.290 ;
        RECT 55.320 48.500 55.950 49.290 ;
        RECT 56.910 48.500 57.540 49.290 ;
        RECT 58.480 48.510 59.110 49.290 ;
        RECT 60.060 48.510 60.690 49.290 ;
        RECT 61.650 48.510 62.280 49.290 ;
        RECT 62.540 49.270 72.070 49.290 ;
        RECT 65.110 48.500 65.740 49.270 ;
        RECT 66.700 48.500 67.330 49.270 ;
        RECT 68.270 48.510 68.900 49.270 ;
        RECT 69.850 48.510 70.480 49.270 ;
        RECT 71.440 48.510 72.070 49.270 ;
        RECT 25.770 38.960 26.400 39.890 ;
        RECT 27.360 38.960 27.990 39.890 ;
        RECT 28.930 38.960 29.560 39.900 ;
        RECT 30.510 38.960 31.140 39.900 ;
        RECT 32.100 38.960 32.730 39.900 ;
        RECT 35.700 38.960 36.330 39.890 ;
        RECT 37.290 38.960 37.920 39.890 ;
        RECT 38.860 38.960 39.490 39.900 ;
        RECT 40.440 38.960 41.070 39.900 ;
        RECT 42.030 38.960 42.660 39.900 ;
        RECT 45.510 38.960 46.140 39.890 ;
        RECT 47.100 38.960 47.730 39.890 ;
        RECT 48.670 38.960 49.300 39.900 ;
        RECT 50.250 38.960 50.880 39.900 ;
        RECT 51.840 38.960 52.470 39.900 ;
        RECT 55.320 38.960 55.950 39.920 ;
        RECT 56.910 38.960 57.540 39.920 ;
        RECT 58.480 38.960 59.110 39.930 ;
        RECT 60.060 38.960 60.690 39.930 ;
        RECT 61.650 38.960 62.280 39.930 ;
        RECT 65.110 38.970 65.740 39.920 ;
        RECT 66.700 38.970 67.330 39.920 ;
        RECT 68.270 38.970 68.900 39.930 ;
        RECT 69.850 38.970 70.480 39.930 ;
        RECT 71.440 38.970 72.070 39.930 ;
        RECT 62.560 38.960 72.070 38.970 ;
        RECT 25.770 36.290 72.070 38.960 ;
        RECT 25.770 35.440 26.400 36.290 ;
        RECT 27.360 35.440 27.990 36.290 ;
        RECT 28.930 35.450 29.560 36.290 ;
        RECT 30.510 35.450 31.140 36.290 ;
        RECT 32.100 35.450 32.730 36.290 ;
        RECT 35.700 35.440 36.330 36.290 ;
        RECT 37.290 35.440 37.920 36.290 ;
        RECT 38.860 35.450 39.490 36.290 ;
        RECT 40.440 35.450 41.070 36.290 ;
        RECT 42.030 35.450 42.660 36.290 ;
        RECT 45.510 35.440 46.140 36.290 ;
        RECT 47.100 35.440 47.730 36.290 ;
        RECT 48.670 35.450 49.300 36.290 ;
        RECT 50.250 35.450 50.880 36.290 ;
        RECT 51.840 35.450 52.470 36.290 ;
        RECT 55.320 35.470 55.950 36.290 ;
        RECT 56.910 35.470 57.540 36.290 ;
        RECT 58.480 35.480 59.110 36.290 ;
        RECT 60.060 35.480 60.690 36.290 ;
        RECT 61.650 35.480 62.280 36.290 ;
        RECT 65.110 35.470 65.740 36.290 ;
        RECT 66.700 35.470 67.330 36.290 ;
        RECT 68.270 35.480 68.900 36.290 ;
        RECT 69.850 35.480 70.480 36.290 ;
        RECT 71.440 35.480 72.070 36.290 ;
        RECT 25.770 27.650 26.400 28.710 ;
        RECT 27.360 27.650 27.990 28.710 ;
        RECT 28.930 27.650 29.560 28.720 ;
        RECT 30.510 27.650 31.140 28.720 ;
        RECT 32.100 27.650 32.730 28.720 ;
        RECT 35.700 27.650 36.330 28.710 ;
        RECT 37.290 27.650 37.920 28.710 ;
        RECT 38.860 27.650 39.490 28.720 ;
        RECT 40.440 27.650 41.070 28.720 ;
        RECT 42.030 27.650 42.660 28.720 ;
        RECT 45.510 27.650 46.140 28.710 ;
        RECT 47.100 27.650 47.730 28.710 ;
        RECT 48.670 27.650 49.300 28.720 ;
        RECT 50.250 27.650 50.880 28.720 ;
        RECT 51.840 27.650 52.470 28.720 ;
        RECT 55.320 27.650 55.950 28.740 ;
        RECT 56.910 27.650 57.540 28.740 ;
        RECT 58.480 27.650 59.110 28.750 ;
        RECT 60.060 27.650 60.690 28.750 ;
        RECT 61.650 27.650 62.280 28.750 ;
        RECT 65.110 27.650 65.740 28.740 ;
        RECT 66.700 27.650 67.330 28.740 ;
        RECT 68.270 27.650 68.900 28.750 ;
        RECT 69.850 27.650 70.480 28.750 ;
        RECT 71.440 27.650 72.070 28.750 ;
        RECT 25.770 24.980 72.070 27.650 ;
        RECT 25.770 24.260 26.400 24.980 ;
        RECT 27.360 24.260 27.990 24.980 ;
        RECT 28.930 24.270 29.560 24.980 ;
        RECT 30.510 24.270 31.140 24.980 ;
        RECT 32.100 24.270 32.730 24.980 ;
        RECT 35.700 24.260 36.330 24.980 ;
        RECT 37.290 24.260 37.920 24.980 ;
        RECT 38.860 24.270 39.490 24.980 ;
        RECT 40.440 24.270 41.070 24.980 ;
        RECT 42.030 24.270 42.660 24.980 ;
        RECT 45.510 24.260 46.140 24.980 ;
        RECT 47.100 24.260 47.730 24.980 ;
        RECT 48.670 24.270 49.300 24.980 ;
        RECT 50.250 24.270 50.880 24.980 ;
        RECT 51.840 24.270 52.470 24.980 ;
        RECT 55.320 24.290 55.950 24.980 ;
        RECT 56.910 24.290 57.540 24.980 ;
        RECT 58.480 24.300 59.110 24.980 ;
        RECT 60.060 24.300 60.690 24.980 ;
        RECT 61.650 24.300 62.280 24.980 ;
        RECT 65.110 24.290 65.740 24.980 ;
        RECT 66.700 24.290 67.330 24.980 ;
        RECT 68.270 24.300 68.900 24.980 ;
        RECT 69.850 24.300 70.480 24.980 ;
        RECT 71.440 24.300 72.070 24.980 ;
        RECT 25.770 16.690 26.400 17.530 ;
        RECT 27.360 16.690 27.990 17.530 ;
        RECT 28.930 16.690 29.560 17.540 ;
        RECT 30.510 16.690 31.140 17.540 ;
        RECT 32.100 16.690 32.730 17.540 ;
        RECT 35.700 16.690 36.330 17.530 ;
        RECT 37.290 16.690 37.920 17.530 ;
        RECT 38.860 16.690 39.490 17.540 ;
        RECT 40.440 16.690 41.070 17.540 ;
        RECT 42.030 16.690 42.660 17.540 ;
        RECT 45.510 16.690 46.140 17.530 ;
        RECT 47.100 16.690 47.730 17.530 ;
        RECT 48.670 16.690 49.300 17.540 ;
        RECT 50.250 16.690 50.880 17.540 ;
        RECT 51.840 16.690 52.470 17.540 ;
        RECT 55.320 16.690 55.950 17.560 ;
        RECT 56.910 16.690 57.540 17.560 ;
        RECT 58.480 16.690 59.110 17.570 ;
        RECT 60.060 16.690 60.690 17.570 ;
        RECT 61.650 16.690 62.280 17.570 ;
        RECT 65.110 16.690 65.740 17.560 ;
        RECT 66.700 16.690 67.330 17.560 ;
        RECT 68.270 16.690 68.900 17.570 ;
        RECT 69.850 16.690 70.480 17.570 ;
        RECT 71.440 16.690 72.070 17.570 ;
        RECT 25.770 14.020 72.070 16.690 ;
        RECT 25.770 13.080 26.400 14.020 ;
        RECT 27.360 13.080 27.990 14.020 ;
        RECT 28.930 13.090 29.560 14.020 ;
        RECT 30.510 13.090 31.140 14.020 ;
        RECT 32.100 13.090 32.730 14.020 ;
        RECT 35.700 13.080 36.330 14.020 ;
        RECT 37.290 13.080 37.920 14.020 ;
        RECT 38.860 13.090 39.490 14.020 ;
        RECT 40.440 13.090 41.070 14.020 ;
        RECT 42.030 13.090 42.660 14.020 ;
        RECT 45.510 13.080 46.140 14.020 ;
        RECT 47.100 13.080 47.730 14.020 ;
        RECT 48.670 13.090 49.300 14.020 ;
        RECT 50.250 13.090 50.880 14.020 ;
        RECT 51.840 13.090 52.470 14.020 ;
        RECT 55.320 13.110 55.950 14.020 ;
        RECT 56.910 13.110 57.540 14.020 ;
        RECT 58.480 13.120 59.110 14.020 ;
        RECT 60.060 13.120 60.690 14.020 ;
        RECT 61.650 13.120 62.280 14.020 ;
        RECT 65.110 13.110 65.740 14.020 ;
        RECT 66.700 13.110 67.330 14.020 ;
        RECT 68.270 13.120 68.900 14.020 ;
        RECT 69.850 13.120 70.480 14.020 ;
        RECT 71.440 13.120 72.070 14.020 ;
        RECT 25.770 5.430 26.400 6.350 ;
        RECT 27.360 5.430 27.990 6.350 ;
        RECT 28.930 5.430 29.560 6.360 ;
        RECT 30.510 5.430 31.140 6.360 ;
        RECT 32.100 5.430 32.730 6.360 ;
        RECT 35.700 5.430 36.330 6.350 ;
        RECT 37.290 5.430 37.920 6.350 ;
        RECT 38.860 5.430 39.490 6.360 ;
        RECT 40.440 5.430 41.070 6.360 ;
        RECT 42.030 5.430 42.660 6.360 ;
        RECT 45.510 5.430 46.140 6.350 ;
        RECT 47.100 5.430 47.730 6.350 ;
        RECT 48.670 5.430 49.300 6.360 ;
        RECT 50.250 5.430 50.880 6.360 ;
        RECT 51.840 5.430 52.470 6.360 ;
        RECT 55.320 5.430 55.950 6.380 ;
        RECT 56.910 5.430 57.540 6.380 ;
        RECT 58.480 5.430 59.110 6.390 ;
        RECT 60.060 5.430 60.690 6.390 ;
        RECT 61.650 5.430 62.280 6.390 ;
        RECT 65.110 5.450 65.740 6.380 ;
        RECT 66.700 5.450 67.330 6.380 ;
        RECT 68.270 5.450 68.900 6.390 ;
        RECT 69.850 5.450 70.480 6.390 ;
        RECT 71.440 5.450 72.070 6.390 ;
        RECT 62.530 5.430 72.070 5.450 ;
        RECT 25.770 2.760 72.070 5.430 ;
        RECT 25.770 1.900 26.400 2.760 ;
        RECT 27.360 1.900 27.990 2.760 ;
        RECT 28.930 1.910 29.560 2.760 ;
        RECT 30.510 1.910 31.140 2.760 ;
        RECT 32.100 1.910 32.730 2.760 ;
        RECT 35.700 1.900 36.330 2.760 ;
        RECT 37.290 1.900 37.920 2.760 ;
        RECT 38.860 1.910 39.490 2.760 ;
        RECT 40.440 1.910 41.070 2.760 ;
        RECT 42.030 1.910 42.660 2.760 ;
        RECT 45.510 1.900 46.140 2.760 ;
        RECT 47.100 1.900 47.730 2.760 ;
        RECT 48.670 1.910 49.300 2.760 ;
        RECT 50.250 1.910 50.880 2.760 ;
        RECT 51.840 1.910 52.470 2.760 ;
        RECT 55.320 1.930 55.950 2.760 ;
        RECT 56.910 1.930 57.540 2.760 ;
        RECT 58.480 1.940 59.110 2.760 ;
        RECT 60.060 1.940 60.690 2.760 ;
        RECT 61.650 1.940 62.280 2.760 ;
        RECT 65.110 1.930 65.740 2.760 ;
        RECT 66.700 1.930 67.330 2.760 ;
        RECT 68.270 1.940 68.900 2.760 ;
        RECT 69.850 1.940 70.480 2.760 ;
        RECT 71.440 1.940 72.070 2.760 ;
      LAYER via2 ;
        RECT 62.530 60.620 71.630 63.170 ;
        RECT 62.540 49.320 71.640 51.870 ;
        RECT 62.560 36.370 71.660 38.920 ;
        RECT 62.530 25.040 71.630 27.590 ;
        RECT 62.530 14.080 71.630 16.630 ;
        RECT 62.530 2.850 71.630 5.400 ;
      LAYER met3 ;
        RECT 62.480 63.050 71.680 63.195 ;
        RECT 62.480 60.595 71.690 63.050 ;
        RECT 62.510 51.895 71.690 60.595 ;
        RECT 62.490 49.295 71.690 51.895 ;
        RECT 62.510 38.945 71.690 49.295 ;
        RECT 62.510 36.345 71.710 38.945 ;
        RECT 62.510 27.615 71.690 36.345 ;
        RECT 62.480 25.015 71.690 27.615 ;
        RECT 62.510 16.655 71.690 25.015 ;
        RECT 62.480 14.055 71.690 16.655 ;
        RECT 62.510 5.425 71.690 14.055 ;
        RECT 62.480 3.000 71.690 5.425 ;
        RECT 62.480 2.825 71.680 3.000 ;
    END
  END out_p
  PIN out_n
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 435.000000 ;
    PORT
      LAYER li1 ;
        RECT 26.030 130.325 26.200 140.365 ;
        RECT 27.610 130.325 27.780 140.365 ;
        RECT 29.190 130.325 29.360 140.365 ;
        RECT 30.770 130.325 30.940 140.365 ;
        RECT 32.350 130.325 32.520 140.365 ;
        RECT 35.970 130.325 36.140 140.365 ;
        RECT 37.550 130.325 37.720 140.365 ;
        RECT 39.130 130.325 39.300 140.365 ;
        RECT 40.710 130.325 40.880 140.365 ;
        RECT 42.290 130.325 42.460 140.365 ;
        RECT 45.770 130.325 45.940 140.365 ;
        RECT 47.350 130.325 47.520 140.365 ;
        RECT 48.930 130.325 49.100 140.365 ;
        RECT 50.510 130.325 50.680 140.365 ;
        RECT 52.090 130.325 52.260 140.365 ;
        RECT 55.570 130.325 55.740 140.365 ;
        RECT 57.150 130.325 57.320 140.365 ;
        RECT 58.730 130.325 58.900 140.365 ;
        RECT 60.310 130.325 60.480 140.365 ;
        RECT 61.890 130.325 62.060 140.365 ;
        RECT 65.370 130.325 65.540 140.365 ;
        RECT 66.950 130.325 67.120 140.365 ;
        RECT 68.530 130.325 68.700 140.365 ;
        RECT 70.110 130.325 70.280 140.365 ;
        RECT 71.690 130.325 71.860 140.365 ;
        RECT 26.030 119.145 26.200 129.185 ;
        RECT 27.610 119.145 27.780 129.185 ;
        RECT 29.190 119.145 29.360 129.185 ;
        RECT 30.770 119.145 30.940 129.185 ;
        RECT 32.350 119.145 32.520 129.185 ;
        RECT 35.970 119.145 36.140 129.185 ;
        RECT 37.550 119.145 37.720 129.185 ;
        RECT 39.130 119.145 39.300 129.185 ;
        RECT 40.710 119.145 40.880 129.185 ;
        RECT 42.290 119.145 42.460 129.185 ;
        RECT 45.770 119.145 45.940 129.185 ;
        RECT 47.350 119.145 47.520 129.185 ;
        RECT 48.930 119.145 49.100 129.185 ;
        RECT 50.510 119.145 50.680 129.185 ;
        RECT 52.090 119.145 52.260 129.185 ;
        RECT 55.570 119.145 55.740 129.185 ;
        RECT 57.150 119.145 57.320 129.185 ;
        RECT 58.730 119.145 58.900 129.185 ;
        RECT 60.310 119.145 60.480 129.185 ;
        RECT 61.890 119.145 62.060 129.185 ;
        RECT 65.370 119.145 65.540 129.185 ;
        RECT 66.950 119.145 67.120 129.185 ;
        RECT 68.530 119.145 68.700 129.185 ;
        RECT 70.110 119.145 70.280 129.185 ;
        RECT 71.690 119.145 71.860 129.185 ;
        RECT 26.030 107.965 26.200 118.005 ;
        RECT 27.610 107.965 27.780 118.005 ;
        RECT 29.190 107.965 29.360 118.005 ;
        RECT 30.770 107.965 30.940 118.005 ;
        RECT 32.350 107.965 32.520 118.005 ;
        RECT 35.970 107.965 36.140 118.005 ;
        RECT 37.550 107.965 37.720 118.005 ;
        RECT 39.130 107.965 39.300 118.005 ;
        RECT 40.710 107.965 40.880 118.005 ;
        RECT 42.290 107.965 42.460 118.005 ;
        RECT 45.770 107.965 45.940 118.005 ;
        RECT 47.350 107.965 47.520 118.005 ;
        RECT 48.930 107.965 49.100 118.005 ;
        RECT 50.510 107.965 50.680 118.005 ;
        RECT 52.090 107.965 52.260 118.005 ;
        RECT 55.570 107.965 55.740 118.005 ;
        RECT 57.150 107.965 57.320 118.005 ;
        RECT 58.730 107.965 58.900 118.005 ;
        RECT 60.310 107.965 60.480 118.005 ;
        RECT 61.890 107.965 62.060 118.005 ;
        RECT 65.370 107.965 65.540 118.005 ;
        RECT 66.950 107.965 67.120 118.005 ;
        RECT 68.530 107.965 68.700 118.005 ;
        RECT 70.110 107.965 70.280 118.005 ;
        RECT 71.690 107.965 71.860 118.005 ;
        RECT 26.030 96.785 26.200 106.825 ;
        RECT 27.610 96.785 27.780 106.825 ;
        RECT 29.190 96.785 29.360 106.825 ;
        RECT 30.770 96.785 30.940 106.825 ;
        RECT 32.350 96.785 32.520 106.825 ;
        RECT 35.970 96.785 36.140 106.825 ;
        RECT 37.550 96.785 37.720 106.825 ;
        RECT 39.130 96.785 39.300 106.825 ;
        RECT 40.710 96.785 40.880 106.825 ;
        RECT 42.290 96.785 42.460 106.825 ;
        RECT 45.770 96.785 45.940 106.825 ;
        RECT 47.350 96.785 47.520 106.825 ;
        RECT 48.930 96.785 49.100 106.825 ;
        RECT 50.510 96.785 50.680 106.825 ;
        RECT 52.090 96.785 52.260 106.825 ;
        RECT 55.570 96.785 55.740 106.825 ;
        RECT 57.150 96.785 57.320 106.825 ;
        RECT 58.730 96.785 58.900 106.825 ;
        RECT 60.310 96.785 60.480 106.825 ;
        RECT 61.890 96.785 62.060 106.825 ;
        RECT 65.370 96.785 65.540 106.825 ;
        RECT 66.950 96.785 67.120 106.825 ;
        RECT 68.530 96.785 68.700 106.825 ;
        RECT 70.110 96.785 70.280 106.825 ;
        RECT 71.690 96.785 71.860 106.825 ;
        RECT 26.035 83.755 26.205 93.795 ;
        RECT 27.615 83.755 27.785 93.795 ;
        RECT 29.195 83.755 29.365 93.795 ;
        RECT 30.775 83.755 30.945 93.795 ;
        RECT 32.355 83.755 32.525 93.795 ;
        RECT 35.975 83.755 36.145 93.795 ;
        RECT 37.555 83.755 37.725 93.795 ;
        RECT 39.135 83.755 39.305 93.795 ;
        RECT 40.715 83.755 40.885 93.795 ;
        RECT 42.295 83.755 42.465 93.795 ;
        RECT 45.775 83.755 45.945 93.795 ;
        RECT 47.355 83.755 47.525 93.795 ;
        RECT 48.935 83.755 49.105 93.795 ;
        RECT 50.515 83.755 50.685 93.795 ;
        RECT 52.095 83.755 52.265 93.795 ;
        RECT 55.575 83.755 55.745 93.795 ;
        RECT 57.155 83.755 57.325 93.795 ;
        RECT 58.735 83.755 58.905 93.795 ;
        RECT 60.315 83.755 60.485 93.795 ;
        RECT 61.895 83.755 62.065 93.795 ;
        RECT 65.375 83.755 65.545 93.795 ;
        RECT 66.955 83.755 67.125 93.795 ;
        RECT 68.535 83.755 68.705 93.795 ;
        RECT 70.115 83.755 70.285 93.795 ;
        RECT 71.695 83.755 71.865 93.795 ;
        RECT 26.035 72.675 26.205 82.715 ;
        RECT 27.615 72.675 27.785 82.715 ;
        RECT 29.195 72.675 29.365 82.715 ;
        RECT 30.775 72.675 30.945 82.715 ;
        RECT 32.355 72.675 32.525 82.715 ;
        RECT 35.975 72.675 36.145 82.715 ;
        RECT 37.555 72.675 37.725 82.715 ;
        RECT 39.135 72.675 39.305 82.715 ;
        RECT 40.715 72.675 40.885 82.715 ;
        RECT 42.295 72.675 42.465 82.715 ;
        RECT 45.775 72.675 45.945 82.715 ;
        RECT 47.355 72.675 47.525 82.715 ;
        RECT 48.935 72.675 49.105 82.715 ;
        RECT 50.515 72.675 50.685 82.715 ;
        RECT 52.095 72.675 52.265 82.715 ;
        RECT 55.575 72.675 55.745 82.715 ;
        RECT 57.155 72.675 57.325 82.715 ;
        RECT 58.735 72.675 58.905 82.715 ;
        RECT 60.315 72.675 60.485 82.715 ;
        RECT 61.895 72.675 62.065 82.715 ;
        RECT 65.375 72.675 65.545 82.715 ;
        RECT 66.955 72.675 67.125 82.715 ;
        RECT 68.535 72.675 68.705 82.715 ;
        RECT 70.115 72.675 70.285 82.715 ;
        RECT 71.695 72.675 71.865 82.715 ;
      LAYER mcon ;
        RECT 26.030 130.405 26.200 140.285 ;
        RECT 27.610 130.405 27.780 140.285 ;
        RECT 29.190 130.405 29.360 140.285 ;
        RECT 30.770 130.405 30.940 140.285 ;
        RECT 32.350 130.405 32.520 140.285 ;
        RECT 35.970 130.405 36.140 140.285 ;
        RECT 37.550 130.405 37.720 140.285 ;
        RECT 39.130 130.405 39.300 140.285 ;
        RECT 40.710 130.405 40.880 140.285 ;
        RECT 42.290 130.405 42.460 140.285 ;
        RECT 45.770 130.405 45.940 140.285 ;
        RECT 47.350 130.405 47.520 140.285 ;
        RECT 48.930 130.405 49.100 140.285 ;
        RECT 50.510 130.405 50.680 140.285 ;
        RECT 52.090 130.405 52.260 140.285 ;
        RECT 55.570 130.405 55.740 140.285 ;
        RECT 57.150 130.405 57.320 140.285 ;
        RECT 58.730 130.405 58.900 140.285 ;
        RECT 60.310 130.405 60.480 140.285 ;
        RECT 61.890 130.405 62.060 140.285 ;
        RECT 65.370 130.405 65.540 140.285 ;
        RECT 66.950 130.405 67.120 140.285 ;
        RECT 68.530 130.405 68.700 140.285 ;
        RECT 70.110 130.405 70.280 140.285 ;
        RECT 71.690 130.405 71.860 140.285 ;
        RECT 26.030 119.225 26.200 129.105 ;
        RECT 27.610 119.225 27.780 129.105 ;
        RECT 29.190 119.225 29.360 129.105 ;
        RECT 30.770 119.225 30.940 129.105 ;
        RECT 32.350 119.225 32.520 129.105 ;
        RECT 35.970 119.225 36.140 129.105 ;
        RECT 37.550 119.225 37.720 129.105 ;
        RECT 39.130 119.225 39.300 129.105 ;
        RECT 40.710 119.225 40.880 129.105 ;
        RECT 42.290 119.225 42.460 129.105 ;
        RECT 45.770 119.225 45.940 129.105 ;
        RECT 47.350 119.225 47.520 129.105 ;
        RECT 48.930 119.225 49.100 129.105 ;
        RECT 50.510 119.225 50.680 129.105 ;
        RECT 52.090 119.225 52.260 129.105 ;
        RECT 55.570 119.225 55.740 129.105 ;
        RECT 57.150 119.225 57.320 129.105 ;
        RECT 58.730 119.225 58.900 129.105 ;
        RECT 60.310 119.225 60.480 129.105 ;
        RECT 61.890 119.225 62.060 129.105 ;
        RECT 65.370 119.225 65.540 129.105 ;
        RECT 66.950 119.225 67.120 129.105 ;
        RECT 68.530 119.225 68.700 129.105 ;
        RECT 70.110 119.225 70.280 129.105 ;
        RECT 71.690 119.225 71.860 129.105 ;
        RECT 26.030 108.045 26.200 117.925 ;
        RECT 27.610 108.045 27.780 117.925 ;
        RECT 29.190 108.045 29.360 117.925 ;
        RECT 30.770 108.045 30.940 117.925 ;
        RECT 32.350 108.045 32.520 117.925 ;
        RECT 35.970 108.045 36.140 117.925 ;
        RECT 37.550 108.045 37.720 117.925 ;
        RECT 39.130 108.045 39.300 117.925 ;
        RECT 40.710 108.045 40.880 117.925 ;
        RECT 42.290 108.045 42.460 117.925 ;
        RECT 45.770 108.045 45.940 117.925 ;
        RECT 47.350 108.045 47.520 117.925 ;
        RECT 48.930 108.045 49.100 117.925 ;
        RECT 50.510 108.045 50.680 117.925 ;
        RECT 52.090 108.045 52.260 117.925 ;
        RECT 55.570 108.045 55.740 117.925 ;
        RECT 57.150 108.045 57.320 117.925 ;
        RECT 58.730 108.045 58.900 117.925 ;
        RECT 60.310 108.045 60.480 117.925 ;
        RECT 61.890 108.045 62.060 117.925 ;
        RECT 65.370 108.045 65.540 117.925 ;
        RECT 66.950 108.045 67.120 117.925 ;
        RECT 68.530 108.045 68.700 117.925 ;
        RECT 70.110 108.045 70.280 117.925 ;
        RECT 71.690 108.045 71.860 117.925 ;
        RECT 26.030 96.865 26.200 106.745 ;
        RECT 27.610 96.865 27.780 106.745 ;
        RECT 29.190 96.865 29.360 106.745 ;
        RECT 30.770 96.865 30.940 106.745 ;
        RECT 32.350 96.865 32.520 106.745 ;
        RECT 35.970 96.865 36.140 106.745 ;
        RECT 37.550 96.865 37.720 106.745 ;
        RECT 39.130 96.865 39.300 106.745 ;
        RECT 40.710 96.865 40.880 106.745 ;
        RECT 42.290 96.865 42.460 106.745 ;
        RECT 45.770 96.865 45.940 106.745 ;
        RECT 47.350 96.865 47.520 106.745 ;
        RECT 48.930 96.865 49.100 106.745 ;
        RECT 50.510 96.865 50.680 106.745 ;
        RECT 52.090 96.865 52.260 106.745 ;
        RECT 55.570 96.865 55.740 106.745 ;
        RECT 57.150 96.865 57.320 106.745 ;
        RECT 58.730 96.865 58.900 106.745 ;
        RECT 60.310 96.865 60.480 106.745 ;
        RECT 61.890 96.865 62.060 106.745 ;
        RECT 65.370 96.865 65.540 106.745 ;
        RECT 66.950 96.865 67.120 106.745 ;
        RECT 68.530 96.865 68.700 106.745 ;
        RECT 70.110 96.865 70.280 106.745 ;
        RECT 71.690 96.865 71.860 106.745 ;
        RECT 26.035 83.835 26.205 93.715 ;
        RECT 27.615 83.835 27.785 93.715 ;
        RECT 29.195 83.835 29.365 93.715 ;
        RECT 30.775 83.835 30.945 93.715 ;
        RECT 32.355 83.835 32.525 93.715 ;
        RECT 35.975 83.835 36.145 93.715 ;
        RECT 37.555 83.835 37.725 93.715 ;
        RECT 39.135 83.835 39.305 93.715 ;
        RECT 40.715 83.835 40.885 93.715 ;
        RECT 42.295 83.835 42.465 93.715 ;
        RECT 45.775 83.835 45.945 93.715 ;
        RECT 47.355 83.835 47.525 93.715 ;
        RECT 48.935 83.835 49.105 93.715 ;
        RECT 50.515 83.835 50.685 93.715 ;
        RECT 52.095 83.835 52.265 93.715 ;
        RECT 55.575 83.835 55.745 93.715 ;
        RECT 57.155 83.835 57.325 93.715 ;
        RECT 58.735 83.835 58.905 93.715 ;
        RECT 60.315 83.835 60.485 93.715 ;
        RECT 61.895 83.835 62.065 93.715 ;
        RECT 65.375 83.835 65.545 93.715 ;
        RECT 66.955 83.835 67.125 93.715 ;
        RECT 68.535 83.835 68.705 93.715 ;
        RECT 70.115 83.835 70.285 93.715 ;
        RECT 71.695 83.835 71.865 93.715 ;
        RECT 26.035 72.755 26.205 82.635 ;
        RECT 27.615 72.755 27.785 82.635 ;
        RECT 29.195 72.755 29.365 82.635 ;
        RECT 30.775 72.755 30.945 82.635 ;
        RECT 32.355 72.755 32.525 82.635 ;
        RECT 35.975 72.755 36.145 82.635 ;
        RECT 37.555 72.755 37.725 82.635 ;
        RECT 39.135 72.755 39.305 82.635 ;
        RECT 40.715 72.755 40.885 82.635 ;
        RECT 42.295 72.755 42.465 82.635 ;
        RECT 45.775 72.755 45.945 82.635 ;
        RECT 47.355 72.755 47.525 82.635 ;
        RECT 48.935 72.755 49.105 82.635 ;
        RECT 50.515 72.755 50.685 82.635 ;
        RECT 52.095 72.755 52.265 82.635 ;
        RECT 55.575 72.755 55.745 82.635 ;
        RECT 57.155 72.755 57.325 82.635 ;
        RECT 58.735 72.755 58.905 82.635 ;
        RECT 60.315 72.755 60.485 82.635 ;
        RECT 61.895 72.755 62.065 82.635 ;
        RECT 65.375 72.755 65.545 82.635 ;
        RECT 66.955 72.755 67.125 82.635 ;
        RECT 68.535 72.755 68.705 82.635 ;
        RECT 70.115 72.755 70.285 82.635 ;
        RECT 71.695 72.755 71.865 82.635 ;
      LAYER met1 ;
        RECT 26.000 139.880 26.230 140.345 ;
        RECT 27.580 139.880 27.810 140.345 ;
        RECT 25.720 135.530 26.450 139.880 ;
        RECT 27.310 135.530 28.040 139.880 ;
        RECT 29.160 139.870 29.390 140.345 ;
        RECT 30.740 139.870 30.970 140.345 ;
        RECT 32.320 139.870 32.550 140.345 ;
        RECT 35.940 139.880 36.170 140.345 ;
        RECT 37.520 139.880 37.750 140.345 ;
        RECT 26.000 130.345 26.230 135.530 ;
        RECT 27.580 130.345 27.810 135.530 ;
        RECT 28.880 135.520 29.610 139.870 ;
        RECT 30.460 135.520 31.190 139.870 ;
        RECT 32.050 135.520 32.780 139.870 ;
        RECT 35.650 135.530 36.380 139.880 ;
        RECT 37.240 135.530 37.970 139.880 ;
        RECT 39.100 139.870 39.330 140.345 ;
        RECT 40.680 139.870 40.910 140.345 ;
        RECT 42.260 139.870 42.490 140.345 ;
        RECT 45.740 139.880 45.970 140.345 ;
        RECT 47.320 139.880 47.550 140.345 ;
        RECT 29.160 130.345 29.390 135.520 ;
        RECT 30.740 130.345 30.970 135.520 ;
        RECT 32.320 130.345 32.550 135.520 ;
        RECT 35.940 130.345 36.170 135.530 ;
        RECT 37.520 130.345 37.750 135.530 ;
        RECT 38.810 135.520 39.540 139.870 ;
        RECT 40.390 135.520 41.120 139.870 ;
        RECT 41.980 135.520 42.710 139.870 ;
        RECT 45.460 135.530 46.190 139.880 ;
        RECT 47.050 135.530 47.780 139.880 ;
        RECT 48.900 139.870 49.130 140.345 ;
        RECT 50.480 139.870 50.710 140.345 ;
        RECT 52.060 139.870 52.290 140.345 ;
        RECT 39.100 130.345 39.330 135.520 ;
        RECT 40.680 130.345 40.910 135.520 ;
        RECT 42.260 130.345 42.490 135.520 ;
        RECT 45.740 130.345 45.970 135.530 ;
        RECT 47.320 130.345 47.550 135.530 ;
        RECT 48.620 135.520 49.350 139.870 ;
        RECT 50.200 135.520 50.930 139.870 ;
        RECT 51.790 135.520 52.520 139.870 ;
        RECT 55.540 139.850 55.770 140.345 ;
        RECT 57.120 139.850 57.350 140.345 ;
        RECT 48.900 130.345 49.130 135.520 ;
        RECT 50.480 130.345 50.710 135.520 ;
        RECT 52.060 130.345 52.290 135.520 ;
        RECT 55.270 135.500 56.000 139.850 ;
        RECT 56.860 135.500 57.590 139.850 ;
        RECT 58.700 139.840 58.930 140.345 ;
        RECT 60.280 139.840 60.510 140.345 ;
        RECT 61.860 139.840 62.090 140.345 ;
        RECT 65.340 139.850 65.570 140.345 ;
        RECT 66.920 139.850 67.150 140.345 ;
        RECT 55.540 130.345 55.770 135.500 ;
        RECT 57.120 130.345 57.350 135.500 ;
        RECT 58.430 135.490 59.160 139.840 ;
        RECT 60.010 135.490 60.740 139.840 ;
        RECT 61.600 135.490 62.330 139.840 ;
        RECT 65.060 135.500 65.790 139.850 ;
        RECT 66.650 135.500 67.380 139.850 ;
        RECT 68.500 139.840 68.730 140.345 ;
        RECT 70.080 139.840 70.310 140.345 ;
        RECT 71.660 139.840 71.890 140.345 ;
        RECT 58.700 130.345 58.930 135.490 ;
        RECT 60.280 130.345 60.510 135.490 ;
        RECT 61.860 130.345 62.090 135.490 ;
        RECT 65.340 130.345 65.570 135.500 ;
        RECT 66.920 130.345 67.150 135.500 ;
        RECT 68.220 135.490 68.950 139.840 ;
        RECT 69.800 135.490 70.530 139.840 ;
        RECT 71.390 135.490 72.120 139.840 ;
        RECT 68.500 130.345 68.730 135.490 ;
        RECT 70.080 130.345 70.310 135.490 ;
        RECT 71.660 130.345 71.890 135.490 ;
        RECT 26.000 128.700 26.230 129.165 ;
        RECT 27.580 128.700 27.810 129.165 ;
        RECT 25.720 124.350 26.450 128.700 ;
        RECT 27.310 124.350 28.040 128.700 ;
        RECT 29.160 128.690 29.390 129.165 ;
        RECT 30.740 128.690 30.970 129.165 ;
        RECT 32.320 128.690 32.550 129.165 ;
        RECT 35.940 128.700 36.170 129.165 ;
        RECT 37.520 128.700 37.750 129.165 ;
        RECT 26.000 119.165 26.230 124.350 ;
        RECT 27.580 119.165 27.810 124.350 ;
        RECT 28.880 124.340 29.610 128.690 ;
        RECT 30.460 124.340 31.190 128.690 ;
        RECT 32.050 124.340 32.780 128.690 ;
        RECT 35.650 124.350 36.380 128.700 ;
        RECT 37.240 124.350 37.970 128.700 ;
        RECT 39.100 128.690 39.330 129.165 ;
        RECT 40.680 128.690 40.910 129.165 ;
        RECT 42.260 128.690 42.490 129.165 ;
        RECT 45.740 128.700 45.970 129.165 ;
        RECT 47.320 128.700 47.550 129.165 ;
        RECT 29.160 119.165 29.390 124.340 ;
        RECT 30.740 119.165 30.970 124.340 ;
        RECT 32.320 119.165 32.550 124.340 ;
        RECT 35.940 119.165 36.170 124.350 ;
        RECT 37.520 119.165 37.750 124.350 ;
        RECT 38.810 124.340 39.540 128.690 ;
        RECT 40.390 124.340 41.120 128.690 ;
        RECT 41.980 124.340 42.710 128.690 ;
        RECT 45.460 124.350 46.190 128.700 ;
        RECT 47.050 124.350 47.780 128.700 ;
        RECT 48.900 128.690 49.130 129.165 ;
        RECT 50.480 128.690 50.710 129.165 ;
        RECT 52.060 128.690 52.290 129.165 ;
        RECT 39.100 119.165 39.330 124.340 ;
        RECT 40.680 119.165 40.910 124.340 ;
        RECT 42.260 119.165 42.490 124.340 ;
        RECT 45.740 119.165 45.970 124.350 ;
        RECT 47.320 119.165 47.550 124.350 ;
        RECT 48.620 124.340 49.350 128.690 ;
        RECT 50.200 124.340 50.930 128.690 ;
        RECT 51.790 124.340 52.520 128.690 ;
        RECT 55.540 128.670 55.770 129.165 ;
        RECT 57.120 128.670 57.350 129.165 ;
        RECT 48.900 119.165 49.130 124.340 ;
        RECT 50.480 119.165 50.710 124.340 ;
        RECT 52.060 119.165 52.290 124.340 ;
        RECT 55.270 124.320 56.000 128.670 ;
        RECT 56.860 124.320 57.590 128.670 ;
        RECT 58.700 128.660 58.930 129.165 ;
        RECT 60.280 128.660 60.510 129.165 ;
        RECT 61.860 128.660 62.090 129.165 ;
        RECT 65.340 128.670 65.570 129.165 ;
        RECT 66.920 128.670 67.150 129.165 ;
        RECT 55.540 119.165 55.770 124.320 ;
        RECT 57.120 119.165 57.350 124.320 ;
        RECT 58.430 124.310 59.160 128.660 ;
        RECT 60.010 124.310 60.740 128.660 ;
        RECT 61.600 124.310 62.330 128.660 ;
        RECT 65.060 124.320 65.790 128.670 ;
        RECT 66.650 124.320 67.380 128.670 ;
        RECT 68.500 128.660 68.730 129.165 ;
        RECT 70.080 128.660 70.310 129.165 ;
        RECT 71.660 128.660 71.890 129.165 ;
        RECT 58.700 119.165 58.930 124.310 ;
        RECT 60.280 119.165 60.510 124.310 ;
        RECT 61.860 119.165 62.090 124.310 ;
        RECT 65.340 119.165 65.570 124.320 ;
        RECT 66.920 119.165 67.150 124.320 ;
        RECT 68.220 124.310 68.950 128.660 ;
        RECT 69.800 124.310 70.530 128.660 ;
        RECT 71.390 124.310 72.120 128.660 ;
        RECT 68.500 119.165 68.730 124.310 ;
        RECT 70.080 119.165 70.310 124.310 ;
        RECT 71.660 119.165 71.890 124.310 ;
        RECT 26.000 117.520 26.230 117.985 ;
        RECT 27.580 117.520 27.810 117.985 ;
        RECT 25.720 113.170 26.450 117.520 ;
        RECT 27.310 113.170 28.040 117.520 ;
        RECT 29.160 117.510 29.390 117.985 ;
        RECT 30.740 117.510 30.970 117.985 ;
        RECT 32.320 117.510 32.550 117.985 ;
        RECT 35.940 117.520 36.170 117.985 ;
        RECT 37.520 117.520 37.750 117.985 ;
        RECT 26.000 107.985 26.230 113.170 ;
        RECT 27.580 107.985 27.810 113.170 ;
        RECT 28.880 113.160 29.610 117.510 ;
        RECT 30.460 113.160 31.190 117.510 ;
        RECT 32.050 113.160 32.780 117.510 ;
        RECT 35.650 113.170 36.380 117.520 ;
        RECT 37.240 113.170 37.970 117.520 ;
        RECT 39.100 117.510 39.330 117.985 ;
        RECT 40.680 117.510 40.910 117.985 ;
        RECT 42.260 117.510 42.490 117.985 ;
        RECT 45.740 117.520 45.970 117.985 ;
        RECT 47.320 117.520 47.550 117.985 ;
        RECT 29.160 107.985 29.390 113.160 ;
        RECT 30.740 107.985 30.970 113.160 ;
        RECT 32.320 107.985 32.550 113.160 ;
        RECT 35.940 107.985 36.170 113.170 ;
        RECT 37.520 107.985 37.750 113.170 ;
        RECT 38.810 113.160 39.540 117.510 ;
        RECT 40.390 113.160 41.120 117.510 ;
        RECT 41.980 113.160 42.710 117.510 ;
        RECT 45.460 113.170 46.190 117.520 ;
        RECT 47.050 113.170 47.780 117.520 ;
        RECT 48.900 117.510 49.130 117.985 ;
        RECT 50.480 117.510 50.710 117.985 ;
        RECT 52.060 117.510 52.290 117.985 ;
        RECT 39.100 107.985 39.330 113.160 ;
        RECT 40.680 107.985 40.910 113.160 ;
        RECT 42.260 107.985 42.490 113.160 ;
        RECT 45.740 107.985 45.970 113.170 ;
        RECT 47.320 107.985 47.550 113.170 ;
        RECT 48.620 113.160 49.350 117.510 ;
        RECT 50.200 113.160 50.930 117.510 ;
        RECT 51.790 113.160 52.520 117.510 ;
        RECT 55.540 117.490 55.770 117.985 ;
        RECT 57.120 117.490 57.350 117.985 ;
        RECT 48.900 107.985 49.130 113.160 ;
        RECT 50.480 107.985 50.710 113.160 ;
        RECT 52.060 107.985 52.290 113.160 ;
        RECT 55.270 113.140 56.000 117.490 ;
        RECT 56.860 113.140 57.590 117.490 ;
        RECT 58.700 117.480 58.930 117.985 ;
        RECT 60.280 117.480 60.510 117.985 ;
        RECT 61.860 117.480 62.090 117.985 ;
        RECT 65.340 117.490 65.570 117.985 ;
        RECT 66.920 117.490 67.150 117.985 ;
        RECT 55.540 107.985 55.770 113.140 ;
        RECT 57.120 107.985 57.350 113.140 ;
        RECT 58.430 113.130 59.160 117.480 ;
        RECT 60.010 113.130 60.740 117.480 ;
        RECT 61.600 113.130 62.330 117.480 ;
        RECT 65.060 113.140 65.790 117.490 ;
        RECT 66.650 113.140 67.380 117.490 ;
        RECT 68.500 117.480 68.730 117.985 ;
        RECT 70.080 117.480 70.310 117.985 ;
        RECT 71.660 117.480 71.890 117.985 ;
        RECT 58.700 107.985 58.930 113.130 ;
        RECT 60.280 107.985 60.510 113.130 ;
        RECT 61.860 107.985 62.090 113.130 ;
        RECT 65.340 107.985 65.570 113.140 ;
        RECT 66.920 107.985 67.150 113.140 ;
        RECT 68.220 113.130 68.950 117.480 ;
        RECT 69.800 113.130 70.530 117.480 ;
        RECT 71.390 113.130 72.120 117.480 ;
        RECT 68.500 107.985 68.730 113.130 ;
        RECT 70.080 107.985 70.310 113.130 ;
        RECT 71.660 107.985 71.890 113.130 ;
        RECT 26.000 106.340 26.230 106.805 ;
        RECT 27.580 106.340 27.810 106.805 ;
        RECT 25.720 101.990 26.450 106.340 ;
        RECT 27.310 101.990 28.040 106.340 ;
        RECT 29.160 106.330 29.390 106.805 ;
        RECT 30.740 106.330 30.970 106.805 ;
        RECT 32.320 106.330 32.550 106.805 ;
        RECT 35.940 106.340 36.170 106.805 ;
        RECT 37.520 106.340 37.750 106.805 ;
        RECT 26.000 96.805 26.230 101.990 ;
        RECT 27.580 96.805 27.810 101.990 ;
        RECT 28.880 101.980 29.610 106.330 ;
        RECT 30.460 101.980 31.190 106.330 ;
        RECT 32.050 101.980 32.780 106.330 ;
        RECT 35.650 101.990 36.380 106.340 ;
        RECT 37.240 101.990 37.970 106.340 ;
        RECT 39.100 106.330 39.330 106.805 ;
        RECT 40.680 106.330 40.910 106.805 ;
        RECT 42.260 106.330 42.490 106.805 ;
        RECT 45.740 106.340 45.970 106.805 ;
        RECT 47.320 106.340 47.550 106.805 ;
        RECT 29.160 96.805 29.390 101.980 ;
        RECT 30.740 96.805 30.970 101.980 ;
        RECT 32.320 96.805 32.550 101.980 ;
        RECT 35.940 96.805 36.170 101.990 ;
        RECT 37.520 96.805 37.750 101.990 ;
        RECT 38.810 101.980 39.540 106.330 ;
        RECT 40.390 101.980 41.120 106.330 ;
        RECT 41.980 101.980 42.710 106.330 ;
        RECT 45.460 101.990 46.190 106.340 ;
        RECT 47.050 101.990 47.780 106.340 ;
        RECT 48.900 106.330 49.130 106.805 ;
        RECT 50.480 106.330 50.710 106.805 ;
        RECT 52.060 106.330 52.290 106.805 ;
        RECT 39.100 96.805 39.330 101.980 ;
        RECT 40.680 96.805 40.910 101.980 ;
        RECT 42.260 96.805 42.490 101.980 ;
        RECT 45.740 96.805 45.970 101.990 ;
        RECT 47.320 96.805 47.550 101.990 ;
        RECT 48.620 101.980 49.350 106.330 ;
        RECT 50.200 101.980 50.930 106.330 ;
        RECT 51.790 101.980 52.520 106.330 ;
        RECT 55.540 106.310 55.770 106.805 ;
        RECT 57.120 106.310 57.350 106.805 ;
        RECT 48.900 96.805 49.130 101.980 ;
        RECT 50.480 96.805 50.710 101.980 ;
        RECT 52.060 96.805 52.290 101.980 ;
        RECT 55.270 101.960 56.000 106.310 ;
        RECT 56.860 101.960 57.590 106.310 ;
        RECT 58.700 106.300 58.930 106.805 ;
        RECT 60.280 106.300 60.510 106.805 ;
        RECT 61.860 106.300 62.090 106.805 ;
        RECT 65.340 106.310 65.570 106.805 ;
        RECT 66.920 106.310 67.150 106.805 ;
        RECT 55.540 96.805 55.770 101.960 ;
        RECT 57.120 96.805 57.350 101.960 ;
        RECT 58.430 101.950 59.160 106.300 ;
        RECT 60.010 101.950 60.740 106.300 ;
        RECT 61.600 101.950 62.330 106.300 ;
        RECT 65.060 101.960 65.790 106.310 ;
        RECT 66.650 101.960 67.380 106.310 ;
        RECT 68.500 106.300 68.730 106.805 ;
        RECT 70.080 106.300 70.310 106.805 ;
        RECT 71.660 106.300 71.890 106.805 ;
        RECT 58.700 96.805 58.930 101.950 ;
        RECT 60.280 96.805 60.510 101.950 ;
        RECT 61.860 96.805 62.090 101.950 ;
        RECT 65.340 96.805 65.570 101.960 ;
        RECT 66.920 96.805 67.150 101.960 ;
        RECT 68.220 101.950 68.950 106.300 ;
        RECT 69.800 101.950 70.530 106.300 ;
        RECT 71.390 101.950 72.120 106.300 ;
        RECT 68.500 96.805 68.730 101.950 ;
        RECT 70.080 96.805 70.310 101.950 ;
        RECT 71.660 96.805 71.890 101.950 ;
        RECT 26.005 93.310 26.235 93.775 ;
        RECT 27.585 93.310 27.815 93.775 ;
        RECT 25.720 88.960 26.450 93.310 ;
        RECT 27.310 88.960 28.040 93.310 ;
        RECT 29.165 93.300 29.395 93.775 ;
        RECT 30.745 93.300 30.975 93.775 ;
        RECT 32.325 93.300 32.555 93.775 ;
        RECT 35.945 93.310 36.175 93.775 ;
        RECT 37.525 93.310 37.755 93.775 ;
        RECT 26.005 83.775 26.235 88.960 ;
        RECT 27.585 83.775 27.815 88.960 ;
        RECT 28.880 88.950 29.610 93.300 ;
        RECT 30.460 88.950 31.190 93.300 ;
        RECT 32.050 88.950 32.780 93.300 ;
        RECT 35.650 88.960 36.380 93.310 ;
        RECT 37.240 88.960 37.970 93.310 ;
        RECT 39.105 93.300 39.335 93.775 ;
        RECT 40.685 93.300 40.915 93.775 ;
        RECT 42.265 93.300 42.495 93.775 ;
        RECT 45.745 93.310 45.975 93.775 ;
        RECT 47.325 93.310 47.555 93.775 ;
        RECT 29.165 83.775 29.395 88.950 ;
        RECT 30.745 83.775 30.975 88.950 ;
        RECT 32.325 83.775 32.555 88.950 ;
        RECT 35.945 83.775 36.175 88.960 ;
        RECT 37.525 83.775 37.755 88.960 ;
        RECT 38.810 88.950 39.540 93.300 ;
        RECT 40.390 88.950 41.120 93.300 ;
        RECT 41.980 88.950 42.710 93.300 ;
        RECT 45.460 88.960 46.190 93.310 ;
        RECT 47.050 88.960 47.780 93.310 ;
        RECT 48.905 93.300 49.135 93.775 ;
        RECT 50.485 93.300 50.715 93.775 ;
        RECT 52.065 93.300 52.295 93.775 ;
        RECT 39.105 83.775 39.335 88.950 ;
        RECT 40.685 83.775 40.915 88.950 ;
        RECT 42.265 83.775 42.495 88.950 ;
        RECT 45.745 83.775 45.975 88.960 ;
        RECT 47.325 83.775 47.555 88.960 ;
        RECT 48.620 88.950 49.350 93.300 ;
        RECT 50.200 88.950 50.930 93.300 ;
        RECT 51.790 88.950 52.520 93.300 ;
        RECT 55.545 93.280 55.775 93.775 ;
        RECT 57.125 93.280 57.355 93.775 ;
        RECT 48.905 83.775 49.135 88.950 ;
        RECT 50.485 83.775 50.715 88.950 ;
        RECT 52.065 83.775 52.295 88.950 ;
        RECT 55.270 88.930 56.000 93.280 ;
        RECT 56.860 88.930 57.590 93.280 ;
        RECT 58.705 93.270 58.935 93.775 ;
        RECT 60.285 93.270 60.515 93.775 ;
        RECT 61.865 93.270 62.095 93.775 ;
        RECT 65.345 93.280 65.575 93.775 ;
        RECT 66.925 93.280 67.155 93.775 ;
        RECT 55.545 83.775 55.775 88.930 ;
        RECT 57.125 83.775 57.355 88.930 ;
        RECT 58.430 88.920 59.160 93.270 ;
        RECT 60.010 88.920 60.740 93.270 ;
        RECT 61.600 88.920 62.330 93.270 ;
        RECT 65.060 88.930 65.790 93.280 ;
        RECT 66.650 88.930 67.380 93.280 ;
        RECT 68.505 93.270 68.735 93.775 ;
        RECT 70.085 93.270 70.315 93.775 ;
        RECT 71.665 93.270 71.895 93.775 ;
        RECT 58.705 83.775 58.935 88.920 ;
        RECT 60.285 83.775 60.515 88.920 ;
        RECT 61.865 83.775 62.095 88.920 ;
        RECT 65.345 83.775 65.575 88.930 ;
        RECT 66.925 83.775 67.155 88.930 ;
        RECT 68.220 88.920 68.950 93.270 ;
        RECT 69.800 88.920 70.530 93.270 ;
        RECT 71.390 88.920 72.120 93.270 ;
        RECT 68.505 83.775 68.735 88.920 ;
        RECT 70.085 83.775 70.315 88.920 ;
        RECT 71.665 83.775 71.895 88.920 ;
        RECT 26.005 82.260 26.235 82.695 ;
        RECT 27.585 82.260 27.815 82.695 ;
        RECT 25.730 77.910 26.460 82.260 ;
        RECT 27.320 77.910 28.050 82.260 ;
        RECT 29.165 82.250 29.395 82.695 ;
        RECT 30.745 82.250 30.975 82.695 ;
        RECT 32.325 82.250 32.555 82.695 ;
        RECT 35.945 82.260 36.175 82.695 ;
        RECT 37.525 82.260 37.755 82.695 ;
        RECT 26.005 72.695 26.235 77.910 ;
        RECT 27.585 72.695 27.815 77.910 ;
        RECT 28.890 77.900 29.620 82.250 ;
        RECT 30.470 77.900 31.200 82.250 ;
        RECT 32.060 77.900 32.790 82.250 ;
        RECT 35.660 77.910 36.390 82.260 ;
        RECT 37.250 77.910 37.980 82.260 ;
        RECT 39.105 82.250 39.335 82.695 ;
        RECT 40.685 82.250 40.915 82.695 ;
        RECT 42.265 82.250 42.495 82.695 ;
        RECT 45.745 82.260 45.975 82.695 ;
        RECT 47.325 82.260 47.555 82.695 ;
        RECT 29.165 72.695 29.395 77.900 ;
        RECT 30.745 72.695 30.975 77.900 ;
        RECT 32.325 72.695 32.555 77.900 ;
        RECT 35.945 72.695 36.175 77.910 ;
        RECT 37.525 72.695 37.755 77.910 ;
        RECT 38.820 77.900 39.550 82.250 ;
        RECT 40.400 77.900 41.130 82.250 ;
        RECT 41.990 77.900 42.720 82.250 ;
        RECT 45.470 77.910 46.200 82.260 ;
        RECT 47.060 77.910 47.790 82.260 ;
        RECT 48.905 82.250 49.135 82.695 ;
        RECT 50.485 82.250 50.715 82.695 ;
        RECT 52.065 82.250 52.295 82.695 ;
        RECT 39.105 72.695 39.335 77.900 ;
        RECT 40.685 72.695 40.915 77.900 ;
        RECT 42.265 72.695 42.495 77.900 ;
        RECT 45.745 72.695 45.975 77.910 ;
        RECT 47.325 72.695 47.555 77.910 ;
        RECT 48.630 77.900 49.360 82.250 ;
        RECT 50.210 77.900 50.940 82.250 ;
        RECT 51.800 77.900 52.530 82.250 ;
        RECT 55.545 82.230 55.775 82.695 ;
        RECT 57.125 82.230 57.355 82.695 ;
        RECT 48.905 72.695 49.135 77.900 ;
        RECT 50.485 72.695 50.715 77.900 ;
        RECT 52.065 72.695 52.295 77.900 ;
        RECT 55.280 77.880 56.010 82.230 ;
        RECT 56.870 77.880 57.600 82.230 ;
        RECT 58.705 82.220 58.935 82.695 ;
        RECT 60.285 82.220 60.515 82.695 ;
        RECT 61.865 82.220 62.095 82.695 ;
        RECT 65.345 82.230 65.575 82.695 ;
        RECT 66.925 82.230 67.155 82.695 ;
        RECT 55.545 72.695 55.775 77.880 ;
        RECT 57.125 72.695 57.355 77.880 ;
        RECT 58.440 77.870 59.170 82.220 ;
        RECT 60.020 77.870 60.750 82.220 ;
        RECT 61.610 77.870 62.340 82.220 ;
        RECT 65.070 77.880 65.800 82.230 ;
        RECT 66.660 77.880 67.390 82.230 ;
        RECT 68.505 82.220 68.735 82.695 ;
        RECT 70.085 82.220 70.315 82.695 ;
        RECT 71.665 82.220 71.895 82.695 ;
        RECT 58.705 72.695 58.935 77.870 ;
        RECT 60.285 72.695 60.515 77.870 ;
        RECT 61.865 72.695 62.095 77.870 ;
        RECT 65.345 72.695 65.575 77.880 ;
        RECT 66.925 72.695 67.155 77.880 ;
        RECT 68.230 77.870 68.960 82.220 ;
        RECT 69.810 77.870 70.540 82.220 ;
        RECT 71.400 77.870 72.130 82.220 ;
        RECT 68.505 72.695 68.735 77.870 ;
        RECT 70.085 72.695 70.315 77.870 ;
        RECT 71.665 72.695 71.895 77.870 ;
      LAYER via ;
        RECT 25.770 135.530 26.400 139.880 ;
        RECT 27.360 135.530 27.990 139.880 ;
        RECT 28.930 135.520 29.560 139.870 ;
        RECT 30.510 135.520 31.140 139.870 ;
        RECT 32.100 135.520 32.730 139.870 ;
        RECT 35.700 135.530 36.330 139.880 ;
        RECT 37.290 135.530 37.920 139.880 ;
        RECT 38.860 135.520 39.490 139.870 ;
        RECT 40.440 135.520 41.070 139.870 ;
        RECT 42.030 135.520 42.660 139.870 ;
        RECT 45.510 135.530 46.140 139.880 ;
        RECT 47.100 135.530 47.730 139.880 ;
        RECT 48.670 135.520 49.300 139.870 ;
        RECT 50.250 135.520 50.880 139.870 ;
        RECT 51.840 135.520 52.470 139.870 ;
        RECT 55.320 135.500 55.950 139.850 ;
        RECT 56.910 135.500 57.540 139.850 ;
        RECT 58.480 135.490 59.110 139.840 ;
        RECT 60.060 135.490 60.690 139.840 ;
        RECT 61.650 135.490 62.280 139.840 ;
        RECT 65.110 135.500 65.740 139.850 ;
        RECT 66.700 135.500 67.330 139.850 ;
        RECT 68.270 135.490 68.900 139.840 ;
        RECT 69.850 135.490 70.480 139.840 ;
        RECT 71.440 135.490 72.070 139.840 ;
        RECT 25.770 124.350 26.400 128.700 ;
        RECT 27.360 124.350 27.990 128.700 ;
        RECT 28.930 124.340 29.560 128.690 ;
        RECT 30.510 124.340 31.140 128.690 ;
        RECT 32.100 124.340 32.730 128.690 ;
        RECT 35.700 124.350 36.330 128.700 ;
        RECT 37.290 124.350 37.920 128.700 ;
        RECT 38.860 124.340 39.490 128.690 ;
        RECT 40.440 124.340 41.070 128.690 ;
        RECT 42.030 124.340 42.660 128.690 ;
        RECT 45.510 124.350 46.140 128.700 ;
        RECT 47.100 124.350 47.730 128.700 ;
        RECT 48.670 124.340 49.300 128.690 ;
        RECT 50.250 124.340 50.880 128.690 ;
        RECT 51.840 124.340 52.470 128.690 ;
        RECT 55.320 124.320 55.950 128.670 ;
        RECT 56.910 124.320 57.540 128.670 ;
        RECT 58.480 124.310 59.110 128.660 ;
        RECT 60.060 124.310 60.690 128.660 ;
        RECT 61.650 124.310 62.280 128.660 ;
        RECT 65.110 124.320 65.740 128.670 ;
        RECT 66.700 124.320 67.330 128.670 ;
        RECT 68.270 124.310 68.900 128.660 ;
        RECT 69.850 124.310 70.480 128.660 ;
        RECT 71.440 124.310 72.070 128.660 ;
        RECT 25.770 113.170 26.400 117.520 ;
        RECT 27.360 113.170 27.990 117.520 ;
        RECT 28.930 113.160 29.560 117.510 ;
        RECT 30.510 113.160 31.140 117.510 ;
        RECT 32.100 113.160 32.730 117.510 ;
        RECT 35.700 113.170 36.330 117.520 ;
        RECT 37.290 113.170 37.920 117.520 ;
        RECT 38.860 113.160 39.490 117.510 ;
        RECT 40.440 113.160 41.070 117.510 ;
        RECT 42.030 113.160 42.660 117.510 ;
        RECT 45.510 113.170 46.140 117.520 ;
        RECT 47.100 113.170 47.730 117.520 ;
        RECT 48.670 113.160 49.300 117.510 ;
        RECT 50.250 113.160 50.880 117.510 ;
        RECT 51.840 113.160 52.470 117.510 ;
        RECT 55.320 113.140 55.950 117.490 ;
        RECT 56.910 113.140 57.540 117.490 ;
        RECT 58.480 113.130 59.110 117.480 ;
        RECT 60.060 113.130 60.690 117.480 ;
        RECT 61.650 113.130 62.280 117.480 ;
        RECT 65.110 113.140 65.740 117.490 ;
        RECT 66.700 113.140 67.330 117.490 ;
        RECT 68.270 113.130 68.900 117.480 ;
        RECT 69.850 113.130 70.480 117.480 ;
        RECT 71.440 113.130 72.070 117.480 ;
        RECT 25.770 101.990 26.400 106.340 ;
        RECT 27.360 101.990 27.990 106.340 ;
        RECT 28.930 101.980 29.560 106.330 ;
        RECT 30.510 101.980 31.140 106.330 ;
        RECT 32.100 101.980 32.730 106.330 ;
        RECT 35.700 101.990 36.330 106.340 ;
        RECT 37.290 101.990 37.920 106.340 ;
        RECT 38.860 101.980 39.490 106.330 ;
        RECT 40.440 101.980 41.070 106.330 ;
        RECT 42.030 101.980 42.660 106.330 ;
        RECT 45.510 101.990 46.140 106.340 ;
        RECT 47.100 101.990 47.730 106.340 ;
        RECT 48.670 101.980 49.300 106.330 ;
        RECT 50.250 101.980 50.880 106.330 ;
        RECT 51.840 101.980 52.470 106.330 ;
        RECT 55.320 101.960 55.950 106.310 ;
        RECT 56.910 101.960 57.540 106.310 ;
        RECT 58.480 101.950 59.110 106.300 ;
        RECT 60.060 101.950 60.690 106.300 ;
        RECT 61.650 101.950 62.280 106.300 ;
        RECT 65.110 101.960 65.740 106.310 ;
        RECT 66.700 101.960 67.330 106.310 ;
        RECT 68.270 101.950 68.900 106.300 ;
        RECT 69.850 101.950 70.480 106.300 ;
        RECT 71.440 101.950 72.070 106.300 ;
        RECT 25.770 88.960 26.400 93.310 ;
        RECT 27.360 88.960 27.990 93.310 ;
        RECT 28.930 88.950 29.560 93.300 ;
        RECT 30.510 88.950 31.140 93.300 ;
        RECT 32.100 88.950 32.730 93.300 ;
        RECT 35.700 88.960 36.330 93.310 ;
        RECT 37.290 88.960 37.920 93.310 ;
        RECT 38.860 88.950 39.490 93.300 ;
        RECT 40.440 88.950 41.070 93.300 ;
        RECT 42.030 88.950 42.660 93.300 ;
        RECT 45.510 88.960 46.140 93.310 ;
        RECT 47.100 88.960 47.730 93.310 ;
        RECT 48.670 88.950 49.300 93.300 ;
        RECT 50.250 88.950 50.880 93.300 ;
        RECT 51.840 88.950 52.470 93.300 ;
        RECT 55.320 88.930 55.950 93.280 ;
        RECT 56.910 88.930 57.540 93.280 ;
        RECT 58.480 88.920 59.110 93.270 ;
        RECT 60.060 88.920 60.690 93.270 ;
        RECT 61.650 88.920 62.280 93.270 ;
        RECT 65.110 88.930 65.740 93.280 ;
        RECT 66.700 88.930 67.330 93.280 ;
        RECT 68.270 88.920 68.900 93.270 ;
        RECT 69.850 88.920 70.480 93.270 ;
        RECT 71.440 88.920 72.070 93.270 ;
        RECT 25.780 77.910 26.410 82.260 ;
        RECT 27.370 77.910 28.000 82.260 ;
        RECT 28.940 77.900 29.570 82.250 ;
        RECT 30.520 77.900 31.150 82.250 ;
        RECT 32.110 77.900 32.740 82.250 ;
        RECT 35.710 77.910 36.340 82.260 ;
        RECT 37.300 77.910 37.930 82.260 ;
        RECT 38.870 77.900 39.500 82.250 ;
        RECT 40.450 77.900 41.080 82.250 ;
        RECT 42.040 77.900 42.670 82.250 ;
        RECT 45.520 77.910 46.150 82.260 ;
        RECT 47.110 77.910 47.740 82.260 ;
        RECT 48.680 77.900 49.310 82.250 ;
        RECT 50.260 77.900 50.890 82.250 ;
        RECT 51.850 77.900 52.480 82.250 ;
        RECT 55.330 77.880 55.960 82.230 ;
        RECT 56.920 77.880 57.550 82.230 ;
        RECT 58.490 77.870 59.120 82.220 ;
        RECT 60.070 77.870 60.700 82.220 ;
        RECT 61.660 77.870 62.290 82.220 ;
        RECT 65.120 77.880 65.750 82.230 ;
        RECT 66.710 77.880 67.340 82.230 ;
        RECT 68.280 77.870 68.910 82.220 ;
        RECT 69.860 77.870 70.490 82.220 ;
        RECT 71.450 77.870 72.080 82.220 ;
      LAYER met2 ;
        RECT 25.770 139.070 26.400 139.930 ;
        RECT 27.360 139.070 27.990 139.930 ;
        RECT 28.930 139.070 29.560 139.920 ;
        RECT 30.510 139.070 31.140 139.920 ;
        RECT 32.100 139.070 32.730 139.920 ;
        RECT 35.700 139.070 36.330 139.930 ;
        RECT 37.290 139.070 37.920 139.930 ;
        RECT 38.860 139.070 39.490 139.920 ;
        RECT 40.440 139.070 41.070 139.920 ;
        RECT 42.030 139.070 42.660 139.920 ;
        RECT 45.510 139.070 46.140 139.930 ;
        RECT 47.100 139.070 47.730 139.930 ;
        RECT 48.670 139.070 49.300 139.920 ;
        RECT 50.250 139.070 50.880 139.920 ;
        RECT 51.840 139.070 52.470 139.920 ;
        RECT 55.320 139.070 55.950 139.900 ;
        RECT 56.910 139.070 57.540 139.900 ;
        RECT 58.480 139.070 59.110 139.890 ;
        RECT 60.060 139.070 60.690 139.890 ;
        RECT 61.650 139.070 62.280 139.890 ;
        RECT 65.110 139.070 65.740 139.900 ;
        RECT 66.700 139.070 67.330 139.900 ;
        RECT 68.270 139.070 68.900 139.890 ;
        RECT 69.850 139.070 70.480 139.890 ;
        RECT 71.440 139.070 72.070 139.890 ;
        RECT 25.770 136.400 72.070 139.070 ;
        RECT 25.770 135.480 26.400 136.400 ;
        RECT 27.360 135.480 27.990 136.400 ;
        RECT 28.930 135.470 29.560 136.400 ;
        RECT 30.510 135.470 31.140 136.400 ;
        RECT 32.100 135.470 32.730 136.400 ;
        RECT 35.700 135.480 36.330 136.400 ;
        RECT 37.290 135.480 37.920 136.400 ;
        RECT 38.860 135.470 39.490 136.400 ;
        RECT 40.440 135.470 41.070 136.400 ;
        RECT 42.030 135.470 42.660 136.400 ;
        RECT 45.510 135.480 46.140 136.400 ;
        RECT 47.100 135.480 47.730 136.400 ;
        RECT 48.670 135.470 49.300 136.400 ;
        RECT 50.250 135.470 50.880 136.400 ;
        RECT 51.840 135.470 52.470 136.400 ;
        RECT 55.320 135.450 55.950 136.400 ;
        RECT 56.910 135.450 57.540 136.400 ;
        RECT 58.480 135.440 59.110 136.400 ;
        RECT 60.060 135.440 60.690 136.400 ;
        RECT 61.650 135.440 62.280 136.400 ;
        RECT 62.530 136.380 72.070 136.400 ;
        RECT 65.110 135.450 65.740 136.380 ;
        RECT 66.700 135.450 67.330 136.380 ;
        RECT 68.270 135.440 68.900 136.380 ;
        RECT 69.850 135.440 70.480 136.380 ;
        RECT 71.440 135.440 72.070 136.380 ;
        RECT 25.770 127.810 26.400 128.750 ;
        RECT 27.360 127.810 27.990 128.750 ;
        RECT 28.930 127.810 29.560 128.740 ;
        RECT 30.510 127.810 31.140 128.740 ;
        RECT 32.100 127.810 32.730 128.740 ;
        RECT 35.700 127.810 36.330 128.750 ;
        RECT 37.290 127.810 37.920 128.750 ;
        RECT 38.860 127.810 39.490 128.740 ;
        RECT 40.440 127.810 41.070 128.740 ;
        RECT 42.030 127.810 42.660 128.740 ;
        RECT 45.510 127.810 46.140 128.750 ;
        RECT 47.100 127.810 47.730 128.750 ;
        RECT 48.670 127.810 49.300 128.740 ;
        RECT 50.250 127.810 50.880 128.740 ;
        RECT 51.840 127.810 52.470 128.740 ;
        RECT 55.320 127.810 55.950 128.720 ;
        RECT 56.910 127.810 57.540 128.720 ;
        RECT 58.480 127.810 59.110 128.710 ;
        RECT 60.060 127.810 60.690 128.710 ;
        RECT 61.650 127.810 62.280 128.710 ;
        RECT 65.110 127.810 65.740 128.720 ;
        RECT 66.700 127.810 67.330 128.720 ;
        RECT 68.270 127.810 68.900 128.710 ;
        RECT 69.850 127.810 70.480 128.710 ;
        RECT 71.440 127.810 72.070 128.710 ;
        RECT 25.770 125.140 72.070 127.810 ;
        RECT 25.770 124.300 26.400 125.140 ;
        RECT 27.360 124.300 27.990 125.140 ;
        RECT 28.930 124.290 29.560 125.140 ;
        RECT 30.510 124.290 31.140 125.140 ;
        RECT 32.100 124.290 32.730 125.140 ;
        RECT 35.700 124.300 36.330 125.140 ;
        RECT 37.290 124.300 37.920 125.140 ;
        RECT 38.860 124.290 39.490 125.140 ;
        RECT 40.440 124.290 41.070 125.140 ;
        RECT 42.030 124.290 42.660 125.140 ;
        RECT 45.510 124.300 46.140 125.140 ;
        RECT 47.100 124.300 47.730 125.140 ;
        RECT 48.670 124.290 49.300 125.140 ;
        RECT 50.250 124.290 50.880 125.140 ;
        RECT 51.840 124.290 52.470 125.140 ;
        RECT 55.320 124.270 55.950 125.140 ;
        RECT 56.910 124.270 57.540 125.140 ;
        RECT 58.480 124.260 59.110 125.140 ;
        RECT 60.060 124.260 60.690 125.140 ;
        RECT 61.650 124.260 62.280 125.140 ;
        RECT 65.110 124.270 65.740 125.140 ;
        RECT 66.700 124.270 67.330 125.140 ;
        RECT 68.270 124.260 68.900 125.140 ;
        RECT 69.850 124.260 70.480 125.140 ;
        RECT 71.440 124.260 72.070 125.140 ;
        RECT 25.770 116.850 26.400 117.570 ;
        RECT 27.360 116.850 27.990 117.570 ;
        RECT 28.930 116.850 29.560 117.560 ;
        RECT 30.510 116.850 31.140 117.560 ;
        RECT 32.100 116.850 32.730 117.560 ;
        RECT 35.700 116.850 36.330 117.570 ;
        RECT 37.290 116.850 37.920 117.570 ;
        RECT 38.860 116.850 39.490 117.560 ;
        RECT 40.440 116.850 41.070 117.560 ;
        RECT 42.030 116.850 42.660 117.560 ;
        RECT 45.510 116.850 46.140 117.570 ;
        RECT 47.100 116.850 47.730 117.570 ;
        RECT 48.670 116.850 49.300 117.560 ;
        RECT 50.250 116.850 50.880 117.560 ;
        RECT 51.840 116.850 52.470 117.560 ;
        RECT 55.320 116.850 55.950 117.540 ;
        RECT 56.910 116.850 57.540 117.540 ;
        RECT 58.480 116.850 59.110 117.530 ;
        RECT 60.060 116.850 60.690 117.530 ;
        RECT 61.650 116.850 62.280 117.530 ;
        RECT 65.110 116.850 65.740 117.540 ;
        RECT 66.700 116.850 67.330 117.540 ;
        RECT 68.270 116.850 68.900 117.530 ;
        RECT 69.850 116.850 70.480 117.530 ;
        RECT 71.440 116.850 72.070 117.530 ;
        RECT 25.770 114.180 72.070 116.850 ;
        RECT 25.770 113.120 26.400 114.180 ;
        RECT 27.360 113.120 27.990 114.180 ;
        RECT 28.930 113.110 29.560 114.180 ;
        RECT 30.510 113.110 31.140 114.180 ;
        RECT 32.100 113.110 32.730 114.180 ;
        RECT 35.700 113.120 36.330 114.180 ;
        RECT 37.290 113.120 37.920 114.180 ;
        RECT 38.860 113.110 39.490 114.180 ;
        RECT 40.440 113.110 41.070 114.180 ;
        RECT 42.030 113.110 42.660 114.180 ;
        RECT 45.510 113.120 46.140 114.180 ;
        RECT 47.100 113.120 47.730 114.180 ;
        RECT 48.670 113.110 49.300 114.180 ;
        RECT 50.250 113.110 50.880 114.180 ;
        RECT 51.840 113.110 52.470 114.180 ;
        RECT 55.320 113.090 55.950 114.180 ;
        RECT 56.910 113.090 57.540 114.180 ;
        RECT 58.480 113.080 59.110 114.180 ;
        RECT 60.060 113.080 60.690 114.180 ;
        RECT 61.650 113.080 62.280 114.180 ;
        RECT 65.110 113.090 65.740 114.180 ;
        RECT 66.700 113.090 67.330 114.180 ;
        RECT 68.270 113.080 68.900 114.180 ;
        RECT 69.850 113.080 70.480 114.180 ;
        RECT 71.440 113.080 72.070 114.180 ;
        RECT 25.770 105.540 26.400 106.390 ;
        RECT 27.360 105.540 27.990 106.390 ;
        RECT 28.930 105.540 29.560 106.380 ;
        RECT 30.510 105.540 31.140 106.380 ;
        RECT 32.100 105.540 32.730 106.380 ;
        RECT 35.700 105.540 36.330 106.390 ;
        RECT 37.290 105.540 37.920 106.390 ;
        RECT 38.860 105.540 39.490 106.380 ;
        RECT 40.440 105.540 41.070 106.380 ;
        RECT 42.030 105.540 42.660 106.380 ;
        RECT 45.510 105.540 46.140 106.390 ;
        RECT 47.100 105.540 47.730 106.390 ;
        RECT 48.670 105.540 49.300 106.380 ;
        RECT 50.250 105.540 50.880 106.380 ;
        RECT 51.840 105.540 52.470 106.380 ;
        RECT 55.320 105.540 55.950 106.360 ;
        RECT 56.910 105.540 57.540 106.360 ;
        RECT 58.480 105.540 59.110 106.350 ;
        RECT 60.060 105.540 60.690 106.350 ;
        RECT 61.650 105.540 62.280 106.350 ;
        RECT 65.110 105.540 65.740 106.360 ;
        RECT 66.700 105.540 67.330 106.360 ;
        RECT 68.270 105.540 68.900 106.350 ;
        RECT 69.850 105.540 70.480 106.350 ;
        RECT 71.440 105.540 72.070 106.350 ;
        RECT 25.770 102.870 72.070 105.540 ;
        RECT 25.770 101.940 26.400 102.870 ;
        RECT 27.360 101.940 27.990 102.870 ;
        RECT 28.930 101.930 29.560 102.870 ;
        RECT 30.510 101.930 31.140 102.870 ;
        RECT 32.100 101.930 32.730 102.870 ;
        RECT 35.700 101.940 36.330 102.870 ;
        RECT 37.290 101.940 37.920 102.870 ;
        RECT 38.860 101.930 39.490 102.870 ;
        RECT 40.440 101.930 41.070 102.870 ;
        RECT 42.030 101.930 42.660 102.870 ;
        RECT 45.510 101.940 46.140 102.870 ;
        RECT 47.100 101.940 47.730 102.870 ;
        RECT 48.670 101.930 49.300 102.870 ;
        RECT 50.250 101.930 50.880 102.870 ;
        RECT 51.840 101.930 52.470 102.870 ;
        RECT 55.320 101.910 55.950 102.870 ;
        RECT 56.910 101.910 57.540 102.870 ;
        RECT 58.480 101.900 59.110 102.870 ;
        RECT 60.060 101.900 60.690 102.870 ;
        RECT 61.650 101.900 62.280 102.870 ;
        RECT 62.560 102.860 72.070 102.870 ;
        RECT 65.110 101.910 65.740 102.860 ;
        RECT 66.700 101.910 67.330 102.860 ;
        RECT 68.270 101.900 68.900 102.860 ;
        RECT 69.850 101.900 70.480 102.860 ;
        RECT 71.440 101.900 72.070 102.860 ;
        RECT 25.770 92.540 26.400 93.360 ;
        RECT 27.360 92.540 27.990 93.360 ;
        RECT 28.930 92.540 29.560 93.350 ;
        RECT 30.510 92.540 31.140 93.350 ;
        RECT 32.100 92.540 32.730 93.350 ;
        RECT 35.700 92.540 36.330 93.360 ;
        RECT 37.290 92.540 37.920 93.360 ;
        RECT 38.860 92.540 39.490 93.350 ;
        RECT 40.440 92.540 41.070 93.350 ;
        RECT 42.030 92.540 42.660 93.350 ;
        RECT 45.510 92.540 46.140 93.360 ;
        RECT 47.100 92.540 47.730 93.360 ;
        RECT 48.670 92.540 49.300 93.350 ;
        RECT 50.250 92.540 50.880 93.350 ;
        RECT 51.840 92.540 52.470 93.350 ;
        RECT 55.320 92.540 55.950 93.330 ;
        RECT 56.910 92.540 57.540 93.330 ;
        RECT 58.480 92.540 59.110 93.320 ;
        RECT 60.060 92.540 60.690 93.320 ;
        RECT 61.650 92.540 62.280 93.320 ;
        RECT 65.110 92.560 65.740 93.330 ;
        RECT 66.700 92.560 67.330 93.330 ;
        RECT 68.270 92.560 68.900 93.320 ;
        RECT 69.850 92.560 70.480 93.320 ;
        RECT 71.440 92.560 72.070 93.320 ;
        RECT 62.540 92.540 72.070 92.560 ;
        RECT 25.770 89.870 72.070 92.540 ;
        RECT 25.770 88.910 26.400 89.870 ;
        RECT 27.360 88.910 27.990 89.870 ;
        RECT 28.930 88.900 29.560 89.870 ;
        RECT 30.510 88.900 31.140 89.870 ;
        RECT 32.100 88.900 32.730 89.870 ;
        RECT 35.700 88.910 36.330 89.870 ;
        RECT 37.290 88.910 37.920 89.870 ;
        RECT 38.860 88.900 39.490 89.870 ;
        RECT 40.440 88.900 41.070 89.870 ;
        RECT 42.030 88.900 42.660 89.870 ;
        RECT 45.510 88.910 46.140 89.870 ;
        RECT 47.100 88.910 47.730 89.870 ;
        RECT 48.670 88.900 49.300 89.870 ;
        RECT 50.250 88.900 50.880 89.870 ;
        RECT 51.840 88.900 52.470 89.870 ;
        RECT 55.320 88.880 55.950 89.870 ;
        RECT 56.910 88.880 57.540 89.870 ;
        RECT 58.480 88.870 59.110 89.870 ;
        RECT 60.060 88.870 60.690 89.870 ;
        RECT 61.650 88.870 62.280 89.870 ;
        RECT 65.110 88.880 65.740 89.870 ;
        RECT 66.700 88.880 67.330 89.870 ;
        RECT 68.270 88.870 68.900 89.870 ;
        RECT 69.850 88.870 70.480 89.870 ;
        RECT 71.440 88.870 72.070 89.870 ;
        RECT 25.780 81.290 26.410 82.310 ;
        RECT 27.370 81.290 28.000 82.310 ;
        RECT 28.940 81.290 29.570 82.300 ;
        RECT 30.520 81.290 31.150 82.300 ;
        RECT 32.110 81.290 32.740 82.300 ;
        RECT 35.710 81.290 36.340 82.310 ;
        RECT 37.300 81.290 37.930 82.310 ;
        RECT 38.870 81.290 39.500 82.300 ;
        RECT 40.450 81.290 41.080 82.300 ;
        RECT 42.040 81.290 42.670 82.300 ;
        RECT 45.520 81.290 46.150 82.310 ;
        RECT 47.110 81.290 47.740 82.310 ;
        RECT 48.680 81.290 49.310 82.300 ;
        RECT 50.260 81.290 50.890 82.300 ;
        RECT 51.850 81.290 52.480 82.300 ;
        RECT 55.330 81.290 55.960 82.280 ;
        RECT 56.920 81.290 57.550 82.280 ;
        RECT 58.490 81.290 59.120 82.270 ;
        RECT 60.070 81.290 60.700 82.270 ;
        RECT 61.660 81.290 62.290 82.270 ;
        RECT 65.120 81.290 65.750 82.280 ;
        RECT 66.710 81.290 67.340 82.280 ;
        RECT 68.280 81.290 68.910 82.270 ;
        RECT 69.860 81.290 70.490 82.270 ;
        RECT 71.450 81.290 72.080 82.270 ;
        RECT 25.780 78.620 72.080 81.290 ;
        RECT 25.780 77.860 26.410 78.620 ;
        RECT 27.370 77.860 28.000 78.620 ;
        RECT 28.940 77.850 29.570 78.620 ;
        RECT 30.520 77.850 31.150 78.620 ;
        RECT 32.110 77.850 32.740 78.620 ;
        RECT 35.710 77.860 36.340 78.620 ;
        RECT 37.300 77.860 37.930 78.620 ;
        RECT 38.870 77.850 39.500 78.620 ;
        RECT 40.450 77.850 41.080 78.620 ;
        RECT 42.040 77.850 42.670 78.620 ;
        RECT 45.520 77.860 46.150 78.620 ;
        RECT 47.110 77.860 47.740 78.620 ;
        RECT 48.680 77.850 49.310 78.620 ;
        RECT 50.260 77.850 50.890 78.620 ;
        RECT 51.850 77.850 52.480 78.620 ;
        RECT 55.330 77.830 55.960 78.620 ;
        RECT 56.920 77.830 57.550 78.620 ;
        RECT 58.490 77.820 59.120 78.620 ;
        RECT 60.070 77.820 60.700 78.620 ;
        RECT 61.660 77.820 62.290 78.620 ;
        RECT 62.530 78.610 72.080 78.620 ;
        RECT 65.120 77.830 65.750 78.610 ;
        RECT 66.710 77.830 67.340 78.610 ;
        RECT 68.280 77.820 68.910 78.610 ;
        RECT 69.860 77.820 70.490 78.610 ;
        RECT 71.450 77.820 72.080 78.610 ;
      LAYER via2 ;
        RECT 62.530 136.430 71.630 138.980 ;
        RECT 62.530 125.200 71.630 127.750 ;
        RECT 62.530 114.240 71.630 116.790 ;
        RECT 62.560 102.910 71.660 105.460 ;
        RECT 62.540 89.960 71.640 92.510 ;
        RECT 62.530 78.660 71.630 81.210 ;
      LAYER met3 ;
        RECT 62.480 138.830 71.680 139.005 ;
        RECT 62.480 136.405 71.690 138.830 ;
        RECT 62.510 127.775 71.690 136.405 ;
        RECT 62.480 125.175 71.690 127.775 ;
        RECT 62.510 116.815 71.690 125.175 ;
        RECT 62.480 114.215 71.690 116.815 ;
        RECT 62.510 105.485 71.690 114.215 ;
        RECT 62.510 102.885 71.710 105.485 ;
        RECT 62.510 92.535 71.690 102.885 ;
        RECT 62.490 89.935 71.690 92.535 ;
        RECT 62.510 81.235 71.690 89.935 ;
        RECT 62.480 78.780 71.690 81.235 ;
        RECT 62.480 78.635 71.680 78.780 ;
    END
  END out_n
  PIN vdd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.340 141.830 12.920 141.930 ;
        RECT 0.340 141.825 14.370 141.830 ;
        RECT 21.460 141.825 73.710 141.830 ;
        RECT 0.340 117.650 73.710 141.825 ;
        RECT 0.340 83.960 12.920 117.650 ;
        RECT 15.250 111.150 73.710 117.650 ;
        RECT 15.245 107.530 73.710 111.150 ;
        RECT 18.735 105.105 73.710 107.530 ;
        RECT 24.170 102.780 73.710 105.105 ;
        RECT 24.180 95.320 73.710 102.780 ;
        RECT 2.305 76.970 13.835 81.930 ;
        RECT 16.675 68.390 23.625 81.360 ;
        RECT 0.240 24.190 12.820 57.970 ;
        RECT 24.180 39.050 73.710 46.510 ;
        RECT 24.170 36.725 73.710 39.050 ;
        RECT 18.735 34.300 73.710 36.725 ;
        RECT 15.245 30.680 73.710 34.300 ;
        RECT 0.240 24.180 13.210 24.190 ;
        RECT 15.250 24.180 73.710 30.680 ;
        RECT 0.240 0.005 73.710 24.180 ;
        RECT 0.240 0.000 14.950 0.005 ;
        RECT 21.460 0.000 73.710 0.005 ;
      LAYER li1 ;
        RECT 0.730 141.370 12.530 141.540 ;
        RECT 23.690 141.435 73.320 141.440 ;
        RECT 0.730 84.520 0.900 141.370 ;
        RECT 1.400 85.425 1.570 140.465 ;
        RECT 11.690 85.425 11.860 140.465 ;
        RECT 12.360 84.520 12.530 141.370 ;
        RECT 14.385 141.265 73.320 141.435 ;
        RECT 14.385 118.245 14.555 141.265 ;
        RECT 23.615 140.970 73.320 141.265 ;
        RECT 15.055 130.325 15.225 140.365 ;
        RECT 16.635 130.325 16.805 140.365 ;
        RECT 18.215 130.325 18.385 140.365 ;
        RECT 19.795 130.325 19.965 140.365 ;
        RECT 21.375 130.325 21.545 140.365 ;
        RECT 22.955 130.325 23.125 140.365 ;
        RECT 15.055 119.145 15.225 129.185 ;
        RECT 16.635 119.145 16.805 129.185 ;
        RECT 18.215 119.145 18.385 129.185 ;
        RECT 19.795 119.145 19.965 129.185 ;
        RECT 21.375 119.145 21.545 129.185 ;
        RECT 22.955 119.145 23.125 129.185 ;
        RECT 23.615 118.245 24.740 140.970 ;
        RECT 25.240 130.325 25.410 140.365 ;
        RECT 26.820 130.325 26.990 140.365 ;
        RECT 28.400 130.325 28.570 140.365 ;
        RECT 29.980 130.325 30.150 140.365 ;
        RECT 31.560 130.325 31.730 140.365 ;
        RECT 33.140 130.325 33.310 140.365 ;
        RECT 25.240 119.145 25.410 129.185 ;
        RECT 26.820 119.145 26.990 129.185 ;
        RECT 28.400 119.145 28.570 129.185 ;
        RECT 29.980 119.145 30.150 129.185 ;
        RECT 31.560 119.145 31.730 129.185 ;
        RECT 33.140 119.145 33.310 129.185 ;
        RECT 14.385 118.075 24.740 118.245 ;
        RECT 15.630 117.570 24.740 118.075 ;
        RECT 15.640 117.505 24.740 117.570 ;
        RECT 15.640 117.500 19.295 117.505 ;
        RECT 15.640 111.660 15.810 117.500 ;
        RECT 16.310 112.560 16.480 116.600 ;
        RECT 17.890 112.560 18.060 116.600 ;
        RECT 18.550 111.660 19.295 117.500 ;
        RECT 15.640 111.590 19.295 111.660 ;
        RECT 15.630 110.640 19.295 111.590 ;
        RECT 15.635 110.590 19.295 110.640 ;
        RECT 15.635 108.090 15.805 110.590 ;
        RECT 17.095 109.000 17.265 110.040 ;
        RECT 18.545 108.090 19.295 110.590 ;
        RECT 15.635 107.920 19.295 108.090 ;
        RECT 19.125 105.665 19.295 107.920 ;
        RECT 19.795 106.565 19.965 116.605 ;
        RECT 21.375 106.565 21.545 116.605 ;
        RECT 22.955 106.565 23.125 116.605 ;
        RECT 23.615 105.665 24.740 117.505 ;
        RECT 25.240 107.965 25.410 118.005 ;
        RECT 26.820 107.965 26.990 118.005 ;
        RECT 28.400 107.965 28.570 118.005 ;
        RECT 29.980 107.965 30.150 118.005 ;
        RECT 31.560 107.965 31.730 118.005 ;
        RECT 33.140 107.965 33.310 118.005 ;
        RECT 19.125 105.495 24.740 105.665 ;
        RECT 23.690 105.480 24.740 105.495 ;
        RECT 24.570 96.160 24.740 105.480 ;
        RECT 25.240 96.785 25.410 106.825 ;
        RECT 26.820 96.785 26.990 106.825 ;
        RECT 28.400 96.785 28.570 106.825 ;
        RECT 29.980 96.785 30.150 106.825 ;
        RECT 31.560 96.785 31.730 106.825 ;
        RECT 33.140 96.785 33.310 106.825 ;
        RECT 33.810 96.160 34.680 140.970 ;
        RECT 35.180 130.325 35.350 140.365 ;
        RECT 36.760 130.325 36.930 140.365 ;
        RECT 38.340 130.325 38.510 140.365 ;
        RECT 39.920 130.325 40.090 140.365 ;
        RECT 41.500 130.325 41.670 140.365 ;
        RECT 43.080 130.325 43.250 140.365 ;
        RECT 35.180 119.145 35.350 129.185 ;
        RECT 36.760 119.145 36.930 129.185 ;
        RECT 38.340 119.145 38.510 129.185 ;
        RECT 39.920 119.145 40.090 129.185 ;
        RECT 41.500 119.145 41.670 129.185 ;
        RECT 43.080 119.145 43.250 129.185 ;
        RECT 35.180 107.965 35.350 118.005 ;
        RECT 36.760 107.965 36.930 118.005 ;
        RECT 38.340 107.965 38.510 118.005 ;
        RECT 39.920 107.965 40.090 118.005 ;
        RECT 41.500 107.965 41.670 118.005 ;
        RECT 43.080 107.965 43.250 118.005 ;
        RECT 35.180 96.785 35.350 106.825 ;
        RECT 36.760 96.785 36.930 106.825 ;
        RECT 38.340 96.785 38.510 106.825 ;
        RECT 39.920 96.785 40.090 106.825 ;
        RECT 41.500 96.785 41.670 106.825 ;
        RECT 43.080 96.785 43.250 106.825 ;
        RECT 43.750 96.160 44.480 140.970 ;
        RECT 44.980 130.325 45.150 140.365 ;
        RECT 46.560 130.325 46.730 140.365 ;
        RECT 48.140 130.325 48.310 140.365 ;
        RECT 49.720 130.325 49.890 140.365 ;
        RECT 51.300 130.325 51.470 140.365 ;
        RECT 52.880 130.325 53.050 140.365 ;
        RECT 44.980 119.145 45.150 129.185 ;
        RECT 46.560 119.145 46.730 129.185 ;
        RECT 48.140 119.145 48.310 129.185 ;
        RECT 49.720 119.145 49.890 129.185 ;
        RECT 51.300 119.145 51.470 129.185 ;
        RECT 52.880 119.145 53.050 129.185 ;
        RECT 44.980 107.965 45.150 118.005 ;
        RECT 46.560 107.965 46.730 118.005 ;
        RECT 48.140 107.965 48.310 118.005 ;
        RECT 49.720 107.965 49.890 118.005 ;
        RECT 51.300 107.965 51.470 118.005 ;
        RECT 52.880 107.965 53.050 118.005 ;
        RECT 44.980 96.785 45.150 106.825 ;
        RECT 46.560 96.785 46.730 106.825 ;
        RECT 48.140 96.785 48.310 106.825 ;
        RECT 49.720 96.785 49.890 106.825 ;
        RECT 51.300 96.785 51.470 106.825 ;
        RECT 52.880 96.785 53.050 106.825 ;
        RECT 53.550 100.410 54.280 140.970 ;
        RECT 54.780 130.325 54.950 140.365 ;
        RECT 56.360 130.325 56.530 140.365 ;
        RECT 57.940 130.325 58.110 140.365 ;
        RECT 59.520 130.325 59.690 140.365 ;
        RECT 61.100 130.325 61.270 140.365 ;
        RECT 62.680 130.325 62.850 140.365 ;
        RECT 54.780 119.145 54.950 129.185 ;
        RECT 56.360 119.145 56.530 129.185 ;
        RECT 57.940 119.145 58.110 129.185 ;
        RECT 59.520 119.145 59.690 129.185 ;
        RECT 61.100 119.145 61.270 129.185 ;
        RECT 62.680 119.145 62.850 129.185 ;
        RECT 54.780 107.965 54.950 118.005 ;
        RECT 56.360 107.965 56.530 118.005 ;
        RECT 57.940 107.965 58.110 118.005 ;
        RECT 59.520 107.965 59.690 118.005 ;
        RECT 61.100 107.965 61.270 118.005 ;
        RECT 62.680 107.965 62.850 118.005 ;
        RECT 53.550 97.990 54.290 100.410 ;
        RECT 53.550 96.160 54.280 97.990 ;
        RECT 54.780 96.785 54.950 106.825 ;
        RECT 56.360 96.785 56.530 106.825 ;
        RECT 57.940 96.785 58.110 106.825 ;
        RECT 59.520 96.785 59.690 106.825 ;
        RECT 61.100 96.785 61.270 106.825 ;
        RECT 62.680 96.785 62.850 106.825 ;
        RECT 63.350 96.160 64.080 140.970 ;
        RECT 64.580 130.325 64.750 140.365 ;
        RECT 66.160 130.325 66.330 140.365 ;
        RECT 67.740 130.325 67.910 140.365 ;
        RECT 69.320 130.325 69.490 140.365 ;
        RECT 70.900 130.325 71.070 140.365 ;
        RECT 72.480 130.325 72.650 140.365 ;
        RECT 64.580 119.145 64.750 129.185 ;
        RECT 66.160 119.145 66.330 129.185 ;
        RECT 67.740 119.145 67.910 129.185 ;
        RECT 69.320 119.145 69.490 129.185 ;
        RECT 70.900 119.145 71.070 129.185 ;
        RECT 72.480 119.145 72.650 129.185 ;
        RECT 64.580 107.965 64.750 118.005 ;
        RECT 66.160 107.965 66.330 118.005 ;
        RECT 67.740 107.965 67.910 118.005 ;
        RECT 69.320 107.965 69.490 118.005 ;
        RECT 70.900 107.965 71.070 118.005 ;
        RECT 72.480 107.965 72.650 118.005 ;
        RECT 64.580 96.785 64.750 106.825 ;
        RECT 66.160 96.785 66.330 106.825 ;
        RECT 67.740 96.785 67.910 106.825 ;
        RECT 69.320 96.785 69.490 106.825 ;
        RECT 70.900 96.785 71.070 106.825 ;
        RECT 72.480 96.785 72.650 106.825 ;
        RECT 73.150 96.160 73.320 140.970 ;
        RECT 24.570 95.710 73.320 96.160 ;
        RECT 0.730 84.350 12.530 84.520 ;
        RECT 2.695 81.370 13.445 81.540 ;
        RECT 2.695 77.530 2.865 81.370 ;
        RECT 3.365 78.430 3.535 80.470 ;
        RECT 4.945 78.430 5.115 80.470 ;
        RECT 6.525 78.430 6.695 80.470 ;
        RECT 7.985 80.455 8.155 81.370 ;
        RECT 7.935 79.855 8.205 80.455 ;
        RECT 7.985 77.530 8.155 79.855 ;
        RECT 9.445 78.430 9.615 80.470 ;
        RECT 11.025 78.430 11.195 80.470 ;
        RECT 12.605 78.430 12.775 80.470 ;
        RECT 13.275 77.530 13.445 81.370 ;
        RECT 2.695 77.360 13.445 77.530 ;
        RECT 17.065 80.800 23.235 80.970 ;
        RECT 17.065 68.950 17.235 80.800 ;
        RECT 17.735 69.850 17.905 79.890 ;
        RECT 19.315 69.850 19.485 79.890 ;
        RECT 19.985 79.800 20.315 80.800 ;
        RECT 19.945 78.950 20.365 79.800 ;
        RECT 19.985 68.950 20.315 78.950 ;
        RECT 20.815 69.850 20.985 79.890 ;
        RECT 22.395 69.850 22.565 79.890 ;
        RECT 23.065 68.950 23.235 80.800 ;
        RECT 17.065 68.780 23.235 68.950 ;
        RECT 0.630 57.410 12.430 57.580 ;
        RECT 0.630 56.500 0.800 57.410 ;
        RECT 12.260 56.510 12.430 57.410 ;
        RECT 1.300 56.500 1.470 56.505 ;
        RECT 0.630 1.460 1.470 56.500 ;
        RECT 11.590 1.460 12.430 56.510 ;
        RECT 24.570 45.670 73.320 46.120 ;
        RECT 24.570 36.350 24.740 45.670 ;
        RECT 23.690 36.335 24.740 36.350 ;
        RECT 19.125 36.165 24.740 36.335 ;
        RECT 19.125 33.910 19.295 36.165 ;
        RECT 15.635 33.740 19.295 33.910 ;
        RECT 15.635 31.240 15.805 33.740 ;
        RECT 17.095 31.790 17.265 32.830 ;
        RECT 18.545 31.240 19.295 33.740 ;
        RECT 15.635 31.190 19.295 31.240 ;
        RECT 15.630 30.240 19.295 31.190 ;
        RECT 15.640 30.170 19.295 30.240 ;
        RECT 15.640 24.330 15.810 30.170 ;
        RECT 16.310 25.230 16.480 29.270 ;
        RECT 17.890 25.230 18.060 29.270 ;
        RECT 18.550 24.330 19.295 30.170 ;
        RECT 19.795 25.225 19.965 35.265 ;
        RECT 21.375 25.225 21.545 35.265 ;
        RECT 22.955 25.225 23.125 35.265 ;
        RECT 15.640 24.325 19.295 24.330 ;
        RECT 23.615 24.325 24.740 36.165 ;
        RECT 25.240 35.005 25.410 45.045 ;
        RECT 26.820 35.005 26.990 45.045 ;
        RECT 28.400 35.005 28.570 45.045 ;
        RECT 29.980 35.005 30.150 45.045 ;
        RECT 31.560 35.005 31.730 45.045 ;
        RECT 33.140 35.005 33.310 45.045 ;
        RECT 15.640 24.260 24.740 24.325 ;
        RECT 15.630 23.755 24.740 24.260 ;
        RECT 25.240 23.825 25.410 33.865 ;
        RECT 26.820 23.825 26.990 33.865 ;
        RECT 28.400 23.825 28.570 33.865 ;
        RECT 29.980 23.825 30.150 33.865 ;
        RECT 31.560 23.825 31.730 33.865 ;
        RECT 33.140 23.825 33.310 33.865 ;
        RECT 0.630 0.560 0.800 1.460 ;
        RECT 12.260 0.560 12.430 1.460 ;
        RECT 0.630 0.390 12.430 0.560 ;
        RECT 14.385 23.585 24.740 23.755 ;
        RECT 14.385 0.565 14.555 23.585 ;
        RECT 15.055 12.645 15.225 22.685 ;
        RECT 16.635 12.645 16.805 22.685 ;
        RECT 18.215 12.645 18.385 22.685 ;
        RECT 19.795 12.645 19.965 22.685 ;
        RECT 21.375 12.645 21.545 22.685 ;
        RECT 22.955 12.645 23.125 22.685 ;
        RECT 15.055 1.465 15.225 11.505 ;
        RECT 16.635 1.465 16.805 11.505 ;
        RECT 18.215 1.465 18.385 11.505 ;
        RECT 19.795 1.465 19.965 11.505 ;
        RECT 21.375 1.465 21.545 11.505 ;
        RECT 22.955 1.465 23.125 11.505 ;
        RECT 23.615 0.860 24.740 23.585 ;
        RECT 25.240 12.645 25.410 22.685 ;
        RECT 26.820 12.645 26.990 22.685 ;
        RECT 28.400 12.645 28.570 22.685 ;
        RECT 29.980 12.645 30.150 22.685 ;
        RECT 31.560 12.645 31.730 22.685 ;
        RECT 33.140 12.645 33.310 22.685 ;
        RECT 25.240 1.465 25.410 11.505 ;
        RECT 26.820 1.465 26.990 11.505 ;
        RECT 28.400 1.465 28.570 11.505 ;
        RECT 29.980 1.465 30.150 11.505 ;
        RECT 31.560 1.465 31.730 11.505 ;
        RECT 33.140 1.465 33.310 11.505 ;
        RECT 33.810 0.860 34.680 45.670 ;
        RECT 35.180 35.005 35.350 45.045 ;
        RECT 36.760 35.005 36.930 45.045 ;
        RECT 38.340 35.005 38.510 45.045 ;
        RECT 39.920 35.005 40.090 45.045 ;
        RECT 41.500 35.005 41.670 45.045 ;
        RECT 43.080 35.005 43.250 45.045 ;
        RECT 35.180 23.825 35.350 33.865 ;
        RECT 36.760 23.825 36.930 33.865 ;
        RECT 38.340 23.825 38.510 33.865 ;
        RECT 39.920 23.825 40.090 33.865 ;
        RECT 41.500 23.825 41.670 33.865 ;
        RECT 43.080 23.825 43.250 33.865 ;
        RECT 35.180 12.645 35.350 22.685 ;
        RECT 36.760 12.645 36.930 22.685 ;
        RECT 38.340 12.645 38.510 22.685 ;
        RECT 39.920 12.645 40.090 22.685 ;
        RECT 41.500 12.645 41.670 22.685 ;
        RECT 43.080 12.645 43.250 22.685 ;
        RECT 35.180 1.465 35.350 11.505 ;
        RECT 36.760 1.465 36.930 11.505 ;
        RECT 38.340 1.465 38.510 11.505 ;
        RECT 39.920 1.465 40.090 11.505 ;
        RECT 41.500 1.465 41.670 11.505 ;
        RECT 43.080 1.465 43.250 11.505 ;
        RECT 43.750 0.860 44.480 45.670 ;
        RECT 44.980 35.005 45.150 45.045 ;
        RECT 46.560 35.005 46.730 45.045 ;
        RECT 48.140 35.005 48.310 45.045 ;
        RECT 49.720 35.005 49.890 45.045 ;
        RECT 51.300 35.005 51.470 45.045 ;
        RECT 52.880 35.005 53.050 45.045 ;
        RECT 53.550 43.840 54.280 45.670 ;
        RECT 53.550 41.420 54.290 43.840 ;
        RECT 44.980 23.825 45.150 33.865 ;
        RECT 46.560 23.825 46.730 33.865 ;
        RECT 48.140 23.825 48.310 33.865 ;
        RECT 49.720 23.825 49.890 33.865 ;
        RECT 51.300 23.825 51.470 33.865 ;
        RECT 52.880 23.825 53.050 33.865 ;
        RECT 44.980 12.645 45.150 22.685 ;
        RECT 46.560 12.645 46.730 22.685 ;
        RECT 48.140 12.645 48.310 22.685 ;
        RECT 49.720 12.645 49.890 22.685 ;
        RECT 51.300 12.645 51.470 22.685 ;
        RECT 52.880 12.645 53.050 22.685 ;
        RECT 44.980 1.465 45.150 11.505 ;
        RECT 46.560 1.465 46.730 11.505 ;
        RECT 48.140 1.465 48.310 11.505 ;
        RECT 49.720 1.465 49.890 11.505 ;
        RECT 51.300 1.465 51.470 11.505 ;
        RECT 52.880 1.465 53.050 11.505 ;
        RECT 53.550 0.860 54.280 41.420 ;
        RECT 54.780 35.005 54.950 45.045 ;
        RECT 56.360 35.005 56.530 45.045 ;
        RECT 57.940 35.005 58.110 45.045 ;
        RECT 59.520 35.005 59.690 45.045 ;
        RECT 61.100 35.005 61.270 45.045 ;
        RECT 62.680 35.005 62.850 45.045 ;
        RECT 54.780 23.825 54.950 33.865 ;
        RECT 56.360 23.825 56.530 33.865 ;
        RECT 57.940 23.825 58.110 33.865 ;
        RECT 59.520 23.825 59.690 33.865 ;
        RECT 61.100 23.825 61.270 33.865 ;
        RECT 62.680 23.825 62.850 33.865 ;
        RECT 54.780 12.645 54.950 22.685 ;
        RECT 56.360 12.645 56.530 22.685 ;
        RECT 57.940 12.645 58.110 22.685 ;
        RECT 59.520 12.645 59.690 22.685 ;
        RECT 61.100 12.645 61.270 22.685 ;
        RECT 62.680 12.645 62.850 22.685 ;
        RECT 54.780 1.465 54.950 11.505 ;
        RECT 56.360 1.465 56.530 11.505 ;
        RECT 57.940 1.465 58.110 11.505 ;
        RECT 59.520 1.465 59.690 11.505 ;
        RECT 61.100 1.465 61.270 11.505 ;
        RECT 62.680 1.465 62.850 11.505 ;
        RECT 63.350 0.860 64.080 45.670 ;
        RECT 64.580 35.005 64.750 45.045 ;
        RECT 66.160 35.005 66.330 45.045 ;
        RECT 67.740 35.005 67.910 45.045 ;
        RECT 69.320 35.005 69.490 45.045 ;
        RECT 70.900 35.005 71.070 45.045 ;
        RECT 72.480 35.005 72.650 45.045 ;
        RECT 64.580 23.825 64.750 33.865 ;
        RECT 66.160 23.825 66.330 33.865 ;
        RECT 67.740 23.825 67.910 33.865 ;
        RECT 69.320 23.825 69.490 33.865 ;
        RECT 70.900 23.825 71.070 33.865 ;
        RECT 72.480 23.825 72.650 33.865 ;
        RECT 64.580 12.645 64.750 22.685 ;
        RECT 66.160 12.645 66.330 22.685 ;
        RECT 67.740 12.645 67.910 22.685 ;
        RECT 69.320 12.645 69.490 22.685 ;
        RECT 70.900 12.645 71.070 22.685 ;
        RECT 72.480 12.645 72.650 22.685 ;
        RECT 64.580 1.465 64.750 11.505 ;
        RECT 66.160 1.465 66.330 11.505 ;
        RECT 67.740 1.465 67.910 11.505 ;
        RECT 69.320 1.465 69.490 11.505 ;
        RECT 70.900 1.465 71.070 11.505 ;
        RECT 72.480 1.465 72.650 11.505 ;
        RECT 73.150 0.860 73.320 45.670 ;
        RECT 23.615 0.565 73.320 0.860 ;
        RECT 14.385 0.395 73.320 0.565 ;
        RECT 23.690 0.390 73.320 0.395 ;
      LAYER mcon ;
        RECT 1.400 85.505 1.570 140.385 ;
        RECT 11.690 85.505 11.860 140.385 ;
        RECT 15.055 130.405 15.225 140.285 ;
        RECT 16.635 130.405 16.805 140.285 ;
        RECT 18.215 130.405 18.385 140.285 ;
        RECT 19.795 130.405 19.965 140.285 ;
        RECT 21.375 130.405 21.545 140.285 ;
        RECT 22.955 130.405 23.125 140.285 ;
        RECT 15.055 119.225 15.225 129.105 ;
        RECT 16.635 119.225 16.805 129.105 ;
        RECT 18.215 119.225 18.385 129.105 ;
        RECT 19.795 119.225 19.965 129.105 ;
        RECT 21.375 119.225 21.545 129.105 ;
        RECT 22.955 119.225 23.125 129.105 ;
        RECT 25.240 130.405 25.410 140.285 ;
        RECT 26.820 130.405 26.990 140.285 ;
        RECT 28.400 130.405 28.570 140.285 ;
        RECT 29.980 130.405 30.150 140.285 ;
        RECT 31.560 130.405 31.730 140.285 ;
        RECT 33.140 130.405 33.310 140.285 ;
        RECT 25.240 119.225 25.410 129.105 ;
        RECT 26.820 119.225 26.990 129.105 ;
        RECT 28.400 119.225 28.570 129.105 ;
        RECT 29.980 119.225 30.150 129.105 ;
        RECT 31.560 119.225 31.730 129.105 ;
        RECT 33.140 119.225 33.310 129.105 ;
        RECT 35.180 130.405 35.350 140.285 ;
        RECT 36.760 130.405 36.930 140.285 ;
        RECT 38.340 130.405 38.510 140.285 ;
        RECT 39.920 130.405 40.090 140.285 ;
        RECT 41.500 130.405 41.670 140.285 ;
        RECT 43.080 130.405 43.250 140.285 ;
        RECT 43.790 131.360 44.480 133.780 ;
        RECT 33.890 120.220 34.580 122.640 ;
        RECT 16.310 112.640 16.480 116.520 ;
        RECT 17.890 112.640 18.060 116.520 ;
        RECT 17.095 109.080 17.265 109.960 ;
        RECT 19.795 106.645 19.965 116.525 ;
        RECT 21.375 106.645 21.545 116.525 ;
        RECT 22.955 106.645 23.125 116.525 ;
        RECT 25.240 108.045 25.410 117.925 ;
        RECT 26.820 108.045 26.990 117.925 ;
        RECT 28.400 108.045 28.570 117.925 ;
        RECT 29.980 108.045 30.150 117.925 ;
        RECT 31.560 108.045 31.730 117.925 ;
        RECT 33.140 108.045 33.310 117.925 ;
        RECT 25.240 96.865 25.410 106.745 ;
        RECT 26.820 96.865 26.990 106.745 ;
        RECT 28.400 96.865 28.570 106.745 ;
        RECT 29.980 96.865 30.150 106.745 ;
        RECT 31.560 96.865 31.730 106.745 ;
        RECT 33.140 96.865 33.310 106.745 ;
        RECT 35.180 119.225 35.350 129.105 ;
        RECT 36.760 119.225 36.930 129.105 ;
        RECT 38.340 119.225 38.510 129.105 ;
        RECT 39.920 119.225 40.090 129.105 ;
        RECT 41.500 119.225 41.670 129.105 ;
        RECT 43.080 119.225 43.250 129.105 ;
        RECT 35.180 108.045 35.350 117.925 ;
        RECT 36.760 108.045 36.930 117.925 ;
        RECT 38.340 108.045 38.510 117.925 ;
        RECT 39.920 108.045 40.090 117.925 ;
        RECT 41.500 108.045 41.670 117.925 ;
        RECT 43.080 108.045 43.250 117.925 ;
        RECT 44.980 130.405 45.150 140.285 ;
        RECT 46.560 130.405 46.730 140.285 ;
        RECT 48.140 130.405 48.310 140.285 ;
        RECT 49.720 130.405 49.890 140.285 ;
        RECT 51.300 130.405 51.470 140.285 ;
        RECT 52.880 130.405 53.050 140.285 ;
        RECT 44.980 119.225 45.150 129.105 ;
        RECT 46.560 119.225 46.730 129.105 ;
        RECT 48.140 119.225 48.310 129.105 ;
        RECT 49.720 119.225 49.890 129.105 ;
        RECT 51.300 119.225 51.470 129.105 ;
        RECT 52.880 119.225 53.050 129.105 ;
        RECT 54.780 130.405 54.950 140.285 ;
        RECT 56.360 130.405 56.530 140.285 ;
        RECT 57.940 130.405 58.110 140.285 ;
        RECT 59.520 130.405 59.690 140.285 ;
        RECT 61.100 130.405 61.270 140.285 ;
        RECT 62.680 130.405 62.850 140.285 ;
        RECT 63.350 131.400 64.040 133.820 ;
        RECT 53.570 120.220 54.260 122.640 ;
        RECT 43.780 108.970 44.470 111.390 ;
        RECT 33.870 98.030 34.560 100.450 ;
        RECT 35.180 96.865 35.350 106.745 ;
        RECT 36.760 96.865 36.930 106.745 ;
        RECT 38.340 96.865 38.510 106.745 ;
        RECT 39.920 96.865 40.090 106.745 ;
        RECT 41.500 96.865 41.670 106.745 ;
        RECT 43.080 96.865 43.250 106.745 ;
        RECT 44.980 108.045 45.150 117.925 ;
        RECT 46.560 108.045 46.730 117.925 ;
        RECT 48.140 108.045 48.310 117.925 ;
        RECT 49.720 108.045 49.890 117.925 ;
        RECT 51.300 108.045 51.470 117.925 ;
        RECT 52.880 108.045 53.050 117.925 ;
        RECT 44.980 96.865 45.150 106.745 ;
        RECT 46.560 96.865 46.730 106.745 ;
        RECT 48.140 96.865 48.310 106.745 ;
        RECT 49.720 96.865 49.890 106.745 ;
        RECT 51.300 96.865 51.470 106.745 ;
        RECT 52.880 96.865 53.050 106.745 ;
        RECT 54.780 119.225 54.950 129.105 ;
        RECT 56.360 119.225 56.530 129.105 ;
        RECT 57.940 119.225 58.110 129.105 ;
        RECT 59.520 119.225 59.690 129.105 ;
        RECT 61.100 119.225 61.270 129.105 ;
        RECT 62.680 119.225 62.850 129.105 ;
        RECT 54.780 108.045 54.950 117.925 ;
        RECT 56.360 108.045 56.530 117.925 ;
        RECT 57.940 108.045 58.110 117.925 ;
        RECT 59.520 108.045 59.690 117.925 ;
        RECT 61.100 108.045 61.270 117.925 ;
        RECT 62.680 108.045 62.850 117.925 ;
        RECT 64.580 130.405 64.750 140.285 ;
        RECT 66.160 130.405 66.330 140.285 ;
        RECT 67.740 130.405 67.910 140.285 ;
        RECT 69.320 130.405 69.490 140.285 ;
        RECT 70.900 130.405 71.070 140.285 ;
        RECT 72.480 130.405 72.650 140.285 ;
        RECT 64.580 119.225 64.750 129.105 ;
        RECT 66.160 119.225 66.330 129.105 ;
        RECT 67.740 119.225 67.910 129.105 ;
        RECT 69.320 119.225 69.490 129.105 ;
        RECT 70.900 119.225 71.070 129.105 ;
        RECT 72.480 119.225 72.650 129.105 ;
        RECT 63.360 108.950 64.050 111.370 ;
        RECT 53.600 97.990 54.290 100.410 ;
        RECT 54.780 96.865 54.950 106.745 ;
        RECT 56.360 96.865 56.530 106.745 ;
        RECT 57.940 96.865 58.110 106.745 ;
        RECT 59.520 96.865 59.690 106.745 ;
        RECT 61.100 96.865 61.270 106.745 ;
        RECT 62.680 96.865 62.850 106.745 ;
        RECT 64.580 108.045 64.750 117.925 ;
        RECT 66.160 108.045 66.330 117.925 ;
        RECT 67.740 108.045 67.910 117.925 ;
        RECT 69.320 108.045 69.490 117.925 ;
        RECT 70.900 108.045 71.070 117.925 ;
        RECT 72.480 108.045 72.650 117.925 ;
        RECT 64.580 96.865 64.750 106.745 ;
        RECT 66.160 96.865 66.330 106.745 ;
        RECT 67.740 96.865 67.910 106.745 ;
        RECT 69.320 96.865 69.490 106.745 ;
        RECT 70.900 96.865 71.070 106.745 ;
        RECT 72.480 96.865 72.650 106.745 ;
        RECT 3.365 78.510 3.535 80.390 ;
        RECT 4.945 78.510 5.115 80.390 ;
        RECT 6.525 78.510 6.695 80.390 ;
        RECT 7.935 79.855 8.205 80.455 ;
        RECT 9.445 78.510 9.615 80.390 ;
        RECT 11.025 78.510 11.195 80.390 ;
        RECT 12.605 78.510 12.775 80.390 ;
        RECT 17.735 69.930 17.905 79.810 ;
        RECT 19.315 69.930 19.485 79.810 ;
        RECT 19.945 78.950 20.365 79.800 ;
        RECT 20.815 69.930 20.985 79.810 ;
        RECT 22.395 69.930 22.565 79.810 ;
        RECT 1.300 1.545 1.470 56.425 ;
        RECT 11.590 1.545 11.760 56.425 ;
        RECT 17.095 31.870 17.265 32.750 ;
        RECT 16.310 25.310 16.480 29.190 ;
        RECT 17.890 25.310 18.060 29.190 ;
        RECT 19.795 25.305 19.965 35.185 ;
        RECT 21.375 25.305 21.545 35.185 ;
        RECT 22.955 25.305 23.125 35.185 ;
        RECT 25.240 35.085 25.410 44.965 ;
        RECT 26.820 35.085 26.990 44.965 ;
        RECT 28.400 35.085 28.570 44.965 ;
        RECT 29.980 35.085 30.150 44.965 ;
        RECT 31.560 35.085 31.730 44.965 ;
        RECT 33.140 35.085 33.310 44.965 ;
        RECT 33.870 41.380 34.560 43.800 ;
        RECT 25.240 23.905 25.410 33.785 ;
        RECT 26.820 23.905 26.990 33.785 ;
        RECT 28.400 23.905 28.570 33.785 ;
        RECT 29.980 23.905 30.150 33.785 ;
        RECT 31.560 23.905 31.730 33.785 ;
        RECT 33.140 23.905 33.310 33.785 ;
        RECT 15.055 12.725 15.225 22.605 ;
        RECT 16.635 12.725 16.805 22.605 ;
        RECT 18.215 12.725 18.385 22.605 ;
        RECT 19.795 12.725 19.965 22.605 ;
        RECT 21.375 12.725 21.545 22.605 ;
        RECT 22.955 12.725 23.125 22.605 ;
        RECT 15.055 1.545 15.225 11.425 ;
        RECT 16.635 1.545 16.805 11.425 ;
        RECT 18.215 1.545 18.385 11.425 ;
        RECT 19.795 1.545 19.965 11.425 ;
        RECT 21.375 1.545 21.545 11.425 ;
        RECT 22.955 1.545 23.125 11.425 ;
        RECT 25.240 12.725 25.410 22.605 ;
        RECT 26.820 12.725 26.990 22.605 ;
        RECT 28.400 12.725 28.570 22.605 ;
        RECT 29.980 12.725 30.150 22.605 ;
        RECT 31.560 12.725 31.730 22.605 ;
        RECT 33.140 12.725 33.310 22.605 ;
        RECT 35.180 35.085 35.350 44.965 ;
        RECT 36.760 35.085 36.930 44.965 ;
        RECT 38.340 35.085 38.510 44.965 ;
        RECT 39.920 35.085 40.090 44.965 ;
        RECT 41.500 35.085 41.670 44.965 ;
        RECT 43.080 35.085 43.250 44.965 ;
        RECT 35.180 23.905 35.350 33.785 ;
        RECT 36.760 23.905 36.930 33.785 ;
        RECT 38.340 23.905 38.510 33.785 ;
        RECT 39.920 23.905 40.090 33.785 ;
        RECT 41.500 23.905 41.670 33.785 ;
        RECT 43.080 23.905 43.250 33.785 ;
        RECT 44.980 35.085 45.150 44.965 ;
        RECT 46.560 35.085 46.730 44.965 ;
        RECT 48.140 35.085 48.310 44.965 ;
        RECT 49.720 35.085 49.890 44.965 ;
        RECT 51.300 35.085 51.470 44.965 ;
        RECT 52.880 35.085 53.050 44.965 ;
        RECT 53.600 41.420 54.290 43.840 ;
        RECT 43.780 30.440 44.470 32.860 ;
        RECT 33.890 19.190 34.580 21.610 ;
        RECT 25.240 1.545 25.410 11.425 ;
        RECT 26.820 1.545 26.990 11.425 ;
        RECT 28.400 1.545 28.570 11.425 ;
        RECT 29.980 1.545 30.150 11.425 ;
        RECT 31.560 1.545 31.730 11.425 ;
        RECT 33.140 1.545 33.310 11.425 ;
        RECT 35.180 12.725 35.350 22.605 ;
        RECT 36.760 12.725 36.930 22.605 ;
        RECT 38.340 12.725 38.510 22.605 ;
        RECT 39.920 12.725 40.090 22.605 ;
        RECT 41.500 12.725 41.670 22.605 ;
        RECT 43.080 12.725 43.250 22.605 ;
        RECT 35.180 1.545 35.350 11.425 ;
        RECT 36.760 1.545 36.930 11.425 ;
        RECT 38.340 1.545 38.510 11.425 ;
        RECT 39.920 1.545 40.090 11.425 ;
        RECT 41.500 1.545 41.670 11.425 ;
        RECT 43.080 1.545 43.250 11.425 ;
        RECT 44.980 23.905 45.150 33.785 ;
        RECT 46.560 23.905 46.730 33.785 ;
        RECT 48.140 23.905 48.310 33.785 ;
        RECT 49.720 23.905 49.890 33.785 ;
        RECT 51.300 23.905 51.470 33.785 ;
        RECT 52.880 23.905 53.050 33.785 ;
        RECT 44.980 12.725 45.150 22.605 ;
        RECT 46.560 12.725 46.730 22.605 ;
        RECT 48.140 12.725 48.310 22.605 ;
        RECT 49.720 12.725 49.890 22.605 ;
        RECT 51.300 12.725 51.470 22.605 ;
        RECT 52.880 12.725 53.050 22.605 ;
        RECT 54.780 35.085 54.950 44.965 ;
        RECT 56.360 35.085 56.530 44.965 ;
        RECT 57.940 35.085 58.110 44.965 ;
        RECT 59.520 35.085 59.690 44.965 ;
        RECT 61.100 35.085 61.270 44.965 ;
        RECT 62.680 35.085 62.850 44.965 ;
        RECT 54.780 23.905 54.950 33.785 ;
        RECT 56.360 23.905 56.530 33.785 ;
        RECT 57.940 23.905 58.110 33.785 ;
        RECT 59.520 23.905 59.690 33.785 ;
        RECT 61.100 23.905 61.270 33.785 ;
        RECT 62.680 23.905 62.850 33.785 ;
        RECT 64.580 35.085 64.750 44.965 ;
        RECT 66.160 35.085 66.330 44.965 ;
        RECT 67.740 35.085 67.910 44.965 ;
        RECT 69.320 35.085 69.490 44.965 ;
        RECT 70.900 35.085 71.070 44.965 ;
        RECT 72.480 35.085 72.650 44.965 ;
        RECT 63.360 30.460 64.050 32.880 ;
        RECT 53.570 19.190 54.260 21.610 ;
        RECT 43.790 8.050 44.480 10.470 ;
        RECT 44.980 1.545 45.150 11.425 ;
        RECT 46.560 1.545 46.730 11.425 ;
        RECT 48.140 1.545 48.310 11.425 ;
        RECT 49.720 1.545 49.890 11.425 ;
        RECT 51.300 1.545 51.470 11.425 ;
        RECT 52.880 1.545 53.050 11.425 ;
        RECT 54.780 12.725 54.950 22.605 ;
        RECT 56.360 12.725 56.530 22.605 ;
        RECT 57.940 12.725 58.110 22.605 ;
        RECT 59.520 12.725 59.690 22.605 ;
        RECT 61.100 12.725 61.270 22.605 ;
        RECT 62.680 12.725 62.850 22.605 ;
        RECT 54.780 1.545 54.950 11.425 ;
        RECT 56.360 1.545 56.530 11.425 ;
        RECT 57.940 1.545 58.110 11.425 ;
        RECT 59.520 1.545 59.690 11.425 ;
        RECT 61.100 1.545 61.270 11.425 ;
        RECT 62.680 1.545 62.850 11.425 ;
        RECT 64.580 23.905 64.750 33.785 ;
        RECT 66.160 23.905 66.330 33.785 ;
        RECT 67.740 23.905 67.910 33.785 ;
        RECT 69.320 23.905 69.490 33.785 ;
        RECT 70.900 23.905 71.070 33.785 ;
        RECT 72.480 23.905 72.650 33.785 ;
        RECT 64.580 12.725 64.750 22.605 ;
        RECT 66.160 12.725 66.330 22.605 ;
        RECT 67.740 12.725 67.910 22.605 ;
        RECT 69.320 12.725 69.490 22.605 ;
        RECT 70.900 12.725 71.070 22.605 ;
        RECT 72.480 12.725 72.650 22.605 ;
        RECT 63.350 8.010 64.040 10.430 ;
        RECT 64.580 1.545 64.750 11.425 ;
        RECT 66.160 1.545 66.330 11.425 ;
        RECT 67.740 1.545 67.910 11.425 ;
        RECT 69.320 1.545 69.490 11.425 ;
        RECT 70.900 1.545 71.070 11.425 ;
        RECT 72.480 1.545 72.650 11.425 ;
      LAYER met1 ;
        RECT 1.370 126.160 1.600 140.445 ;
        RECT 11.660 126.160 11.890 140.445 ;
        RECT 15.025 139.870 15.255 140.345 ;
        RECT 16.605 139.880 16.835 140.345 ;
        RECT 14.950 139.220 15.350 139.870 ;
        RECT 16.510 139.230 16.910 139.880 ;
        RECT 18.185 139.870 18.415 140.345 ;
        RECT 19.765 139.880 19.995 140.345 ;
        RECT 15.025 130.345 15.255 139.220 ;
        RECT 16.605 130.345 16.835 139.230 ;
        RECT 18.110 139.220 18.510 139.870 ;
        RECT 19.680 139.230 20.080 139.880 ;
        RECT 21.345 139.870 21.575 140.345 ;
        RECT 22.925 139.870 23.155 140.345 ;
        RECT 18.185 130.345 18.415 139.220 ;
        RECT 19.765 130.345 19.995 139.230 ;
        RECT 21.260 139.220 21.660 139.870 ;
        RECT 22.840 139.220 23.240 139.870 ;
        RECT 21.345 130.345 21.575 139.220 ;
        RECT 22.925 130.345 23.155 139.220 ;
        RECT 25.210 134.940 25.440 140.345 ;
        RECT 26.790 134.940 27.020 140.345 ;
        RECT 24.950 130.590 25.680 134.940 ;
        RECT 26.540 130.590 27.270 134.940 ;
        RECT 28.370 134.930 28.600 140.345 ;
        RECT 29.950 134.930 30.180 140.345 ;
        RECT 31.530 134.930 31.760 140.345 ;
        RECT 33.110 134.930 33.340 140.345 ;
        RECT 35.150 134.940 35.380 140.345 ;
        RECT 36.730 134.940 36.960 140.345 ;
        RECT 25.210 130.345 25.440 130.590 ;
        RECT 26.790 130.345 27.020 130.590 ;
        RECT 28.110 130.580 28.840 134.930 ;
        RECT 29.690 130.580 30.420 134.930 ;
        RECT 31.280 130.580 32.010 134.930 ;
        RECT 32.850 130.580 33.580 134.930 ;
        RECT 34.880 130.590 35.610 134.940 ;
        RECT 36.470 130.590 37.200 134.940 ;
        RECT 38.310 134.930 38.540 140.345 ;
        RECT 39.890 134.930 40.120 140.345 ;
        RECT 41.470 134.930 41.700 140.345 ;
        RECT 43.050 134.930 43.280 140.345 ;
        RECT 44.950 134.940 45.180 140.345 ;
        RECT 46.530 134.940 46.760 140.345 ;
        RECT 28.370 130.345 28.600 130.580 ;
        RECT 29.950 130.345 30.180 130.580 ;
        RECT 31.530 130.345 31.760 130.580 ;
        RECT 33.110 130.345 33.340 130.580 ;
        RECT 35.150 130.345 35.380 130.590 ;
        RECT 36.730 130.345 36.960 130.590 ;
        RECT 38.040 130.580 38.770 134.930 ;
        RECT 39.620 130.580 40.350 134.930 ;
        RECT 41.210 130.580 41.940 134.930 ;
        RECT 42.780 130.580 43.510 134.930 ;
        RECT 43.760 133.780 44.510 133.840 ;
        RECT 43.740 131.360 44.530 133.780 ;
        RECT 43.760 131.300 44.510 131.360 ;
        RECT 44.690 130.590 45.420 134.940 ;
        RECT 46.280 130.590 47.010 134.940 ;
        RECT 48.110 134.930 48.340 140.345 ;
        RECT 49.690 134.930 49.920 140.345 ;
        RECT 51.270 134.930 51.500 140.345 ;
        RECT 52.850 134.930 53.080 140.345 ;
        RECT 38.310 130.345 38.540 130.580 ;
        RECT 39.890 130.345 40.120 130.580 ;
        RECT 41.470 130.345 41.700 130.580 ;
        RECT 43.050 130.345 43.280 130.580 ;
        RECT 44.950 130.345 45.180 130.590 ;
        RECT 46.530 130.345 46.760 130.590 ;
        RECT 47.850 130.580 48.580 134.930 ;
        RECT 49.430 130.580 50.160 134.930 ;
        RECT 51.020 130.580 51.750 134.930 ;
        RECT 52.590 130.580 53.320 134.930 ;
        RECT 54.750 134.910 54.980 140.345 ;
        RECT 56.330 134.910 56.560 140.345 ;
        RECT 48.110 130.345 48.340 130.580 ;
        RECT 49.690 130.345 49.920 130.580 ;
        RECT 51.270 130.345 51.500 130.580 ;
        RECT 52.850 130.345 53.080 130.580 ;
        RECT 54.500 130.560 55.230 134.910 ;
        RECT 56.090 130.560 56.820 134.910 ;
        RECT 57.910 134.900 58.140 140.345 ;
        RECT 59.490 134.900 59.720 140.345 ;
        RECT 61.070 134.900 61.300 140.345 ;
        RECT 62.650 134.900 62.880 140.345 ;
        RECT 64.550 134.910 64.780 140.345 ;
        RECT 66.130 134.910 66.360 140.345 ;
        RECT 54.750 130.345 54.980 130.560 ;
        RECT 56.330 130.345 56.560 130.560 ;
        RECT 57.660 130.550 58.390 134.900 ;
        RECT 59.240 130.550 59.970 134.900 ;
        RECT 60.830 130.550 61.560 134.900 ;
        RECT 62.400 130.550 63.130 134.900 ;
        RECT 63.320 133.820 64.070 133.880 ;
        RECT 63.300 131.400 64.090 133.820 ;
        RECT 63.320 131.340 64.070 131.400 ;
        RECT 64.290 130.560 65.020 134.910 ;
        RECT 65.880 130.560 66.610 134.910 ;
        RECT 67.710 134.900 67.940 140.345 ;
        RECT 69.290 134.900 69.520 140.345 ;
        RECT 70.870 134.900 71.100 140.345 ;
        RECT 72.450 134.900 72.680 140.345 ;
        RECT 57.910 130.345 58.140 130.550 ;
        RECT 59.490 130.345 59.720 130.550 ;
        RECT 61.070 130.345 61.300 130.550 ;
        RECT 62.650 130.345 62.880 130.550 ;
        RECT 64.550 130.345 64.780 130.560 ;
        RECT 66.130 130.345 66.360 130.560 ;
        RECT 67.450 130.550 68.180 134.900 ;
        RECT 69.030 130.550 69.760 134.900 ;
        RECT 70.620 130.550 71.350 134.900 ;
        RECT 72.190 130.550 72.920 134.900 ;
        RECT 67.710 130.345 67.940 130.550 ;
        RECT 69.290 130.345 69.520 130.550 ;
        RECT 70.870 130.345 71.100 130.550 ;
        RECT 72.450 130.345 72.680 130.550 ;
        RECT 1.370 116.030 11.890 126.160 ;
        RECT 15.025 120.470 15.255 129.165 ;
        RECT 16.605 120.480 16.835 129.165 ;
        RECT 14.930 119.820 15.330 120.470 ;
        RECT 16.510 119.830 16.910 120.480 ;
        RECT 18.185 120.470 18.415 129.165 ;
        RECT 15.025 119.165 15.255 119.820 ;
        RECT 16.605 119.165 16.835 119.830 ;
        RECT 18.080 119.820 18.480 120.470 ;
        RECT 19.765 120.460 19.995 129.165 ;
        RECT 21.345 120.460 21.575 129.165 ;
        RECT 22.925 120.460 23.155 129.165 ;
        RECT 25.210 123.760 25.440 129.165 ;
        RECT 26.790 123.760 27.020 129.165 ;
        RECT 18.185 119.165 18.415 119.820 ;
        RECT 19.680 119.810 20.080 120.460 ;
        RECT 21.260 119.810 21.660 120.460 ;
        RECT 22.840 119.810 23.240 120.460 ;
        RECT 19.765 119.165 19.995 119.810 ;
        RECT 21.345 119.165 21.575 119.810 ;
        RECT 22.925 119.165 23.155 119.810 ;
        RECT 24.950 119.410 25.680 123.760 ;
        RECT 26.540 119.410 27.270 123.760 ;
        RECT 28.370 123.750 28.600 129.165 ;
        RECT 29.950 123.750 30.180 129.165 ;
        RECT 31.530 123.750 31.760 129.165 ;
        RECT 33.110 123.750 33.340 129.165 ;
        RECT 35.150 123.760 35.380 129.165 ;
        RECT 36.730 123.760 36.960 129.165 ;
        RECT 25.210 119.165 25.440 119.410 ;
        RECT 26.790 119.165 27.020 119.410 ;
        RECT 28.110 119.400 28.840 123.750 ;
        RECT 29.690 119.400 30.420 123.750 ;
        RECT 31.280 119.400 32.010 123.750 ;
        RECT 32.850 119.400 33.580 123.750 ;
        RECT 33.860 122.640 34.610 122.700 ;
        RECT 33.840 120.220 34.630 122.640 ;
        RECT 33.860 120.160 34.610 120.220 ;
        RECT 34.880 119.410 35.610 123.760 ;
        RECT 36.470 119.410 37.200 123.760 ;
        RECT 38.310 123.750 38.540 129.165 ;
        RECT 39.890 123.750 40.120 129.165 ;
        RECT 41.470 123.750 41.700 129.165 ;
        RECT 43.050 123.750 43.280 129.165 ;
        RECT 44.950 123.760 45.180 129.165 ;
        RECT 46.530 123.760 46.760 129.165 ;
        RECT 28.370 119.165 28.600 119.400 ;
        RECT 29.950 119.165 30.180 119.400 ;
        RECT 31.530 119.165 31.760 119.400 ;
        RECT 33.110 119.165 33.340 119.400 ;
        RECT 35.150 119.165 35.380 119.410 ;
        RECT 36.730 119.165 36.960 119.410 ;
        RECT 38.040 119.400 38.770 123.750 ;
        RECT 39.620 119.400 40.350 123.750 ;
        RECT 41.210 119.400 41.940 123.750 ;
        RECT 42.780 119.400 43.510 123.750 ;
        RECT 44.690 119.410 45.420 123.760 ;
        RECT 46.280 119.410 47.010 123.760 ;
        RECT 48.110 123.750 48.340 129.165 ;
        RECT 49.690 123.750 49.920 129.165 ;
        RECT 51.270 123.750 51.500 129.165 ;
        RECT 52.850 123.750 53.080 129.165 ;
        RECT 38.310 119.165 38.540 119.400 ;
        RECT 39.890 119.165 40.120 119.400 ;
        RECT 41.470 119.165 41.700 119.400 ;
        RECT 43.050 119.165 43.280 119.400 ;
        RECT 44.950 119.165 45.180 119.410 ;
        RECT 46.530 119.165 46.760 119.410 ;
        RECT 47.850 119.400 48.580 123.750 ;
        RECT 49.430 119.400 50.160 123.750 ;
        RECT 51.020 119.400 51.750 123.750 ;
        RECT 52.590 119.400 53.320 123.750 ;
        RECT 54.750 123.730 54.980 129.165 ;
        RECT 56.330 123.730 56.560 129.165 ;
        RECT 53.540 122.640 54.290 122.700 ;
        RECT 53.520 120.220 54.310 122.640 ;
        RECT 53.540 120.160 54.290 120.220 ;
        RECT 48.110 119.165 48.340 119.400 ;
        RECT 49.690 119.165 49.920 119.400 ;
        RECT 51.270 119.165 51.500 119.400 ;
        RECT 52.850 119.165 53.080 119.400 ;
        RECT 54.500 119.380 55.230 123.730 ;
        RECT 56.090 119.380 56.820 123.730 ;
        RECT 57.910 123.720 58.140 129.165 ;
        RECT 59.490 123.720 59.720 129.165 ;
        RECT 61.070 123.720 61.300 129.165 ;
        RECT 62.650 123.720 62.880 129.165 ;
        RECT 64.550 123.730 64.780 129.165 ;
        RECT 66.130 123.730 66.360 129.165 ;
        RECT 54.750 119.165 54.980 119.380 ;
        RECT 56.330 119.165 56.560 119.380 ;
        RECT 57.660 119.370 58.390 123.720 ;
        RECT 59.240 119.370 59.970 123.720 ;
        RECT 60.830 119.370 61.560 123.720 ;
        RECT 62.400 119.370 63.130 123.720 ;
        RECT 64.290 119.380 65.020 123.730 ;
        RECT 65.880 119.380 66.610 123.730 ;
        RECT 67.710 123.720 67.940 129.165 ;
        RECT 69.290 123.720 69.520 129.165 ;
        RECT 70.870 123.720 71.100 129.165 ;
        RECT 72.450 123.720 72.680 129.165 ;
        RECT 57.910 119.165 58.140 119.370 ;
        RECT 59.490 119.165 59.720 119.370 ;
        RECT 61.070 119.165 61.300 119.370 ;
        RECT 62.650 119.165 62.880 119.370 ;
        RECT 64.550 119.165 64.780 119.380 ;
        RECT 66.130 119.165 66.360 119.380 ;
        RECT 67.450 119.370 68.180 123.720 ;
        RECT 69.030 119.370 69.760 123.720 ;
        RECT 70.620 119.370 71.350 123.720 ;
        RECT 72.190 119.370 72.920 123.720 ;
        RECT 67.710 119.165 67.940 119.370 ;
        RECT 69.290 119.165 69.520 119.370 ;
        RECT 70.870 119.165 71.100 119.370 ;
        RECT 72.450 119.165 72.680 119.370 ;
        RECT 1.370 85.445 1.600 116.030 ;
        RECT 11.660 85.445 11.890 116.030 ;
        RECT 16.280 115.960 16.510 116.580 ;
        RECT 17.860 115.960 18.090 116.580 ;
        RECT 19.765 116.000 19.995 116.585 ;
        RECT 16.200 115.310 16.600 115.960 ;
        RECT 17.760 115.310 18.160 115.960 ;
        RECT 19.670 115.350 20.070 116.000 ;
        RECT 21.345 115.970 21.575 116.585 ;
        RECT 22.925 115.970 23.155 116.585 ;
        RECT 16.280 112.580 16.510 115.310 ;
        RECT 17.860 112.580 18.090 115.310 ;
        RECT 17.065 109.870 17.295 110.020 ;
        RECT 16.980 109.220 17.380 109.870 ;
        RECT 17.065 109.020 17.295 109.220 ;
        RECT 19.765 106.585 19.995 115.350 ;
        RECT 21.260 115.320 21.660 115.970 ;
        RECT 22.820 115.320 23.220 115.970 ;
        RECT 21.345 106.585 21.575 115.320 ;
        RECT 22.925 106.585 23.155 115.320 ;
        RECT 25.210 112.580 25.440 117.985 ;
        RECT 26.790 112.580 27.020 117.985 ;
        RECT 24.950 108.230 25.680 112.580 ;
        RECT 26.540 108.230 27.270 112.580 ;
        RECT 28.370 112.570 28.600 117.985 ;
        RECT 29.950 112.570 30.180 117.985 ;
        RECT 31.530 112.570 31.760 117.985 ;
        RECT 33.110 112.570 33.340 117.985 ;
        RECT 35.150 112.580 35.380 117.985 ;
        RECT 36.730 112.580 36.960 117.985 ;
        RECT 25.210 107.985 25.440 108.230 ;
        RECT 26.790 107.985 27.020 108.230 ;
        RECT 28.110 108.220 28.840 112.570 ;
        RECT 29.690 108.220 30.420 112.570 ;
        RECT 31.280 108.220 32.010 112.570 ;
        RECT 32.850 108.220 33.580 112.570 ;
        RECT 34.880 108.230 35.610 112.580 ;
        RECT 36.470 108.230 37.200 112.580 ;
        RECT 38.310 112.570 38.540 117.985 ;
        RECT 39.890 112.570 40.120 117.985 ;
        RECT 41.470 112.570 41.700 117.985 ;
        RECT 43.050 112.570 43.280 117.985 ;
        RECT 44.950 112.580 45.180 117.985 ;
        RECT 46.530 112.580 46.760 117.985 ;
        RECT 28.370 107.985 28.600 108.220 ;
        RECT 29.950 107.985 30.180 108.220 ;
        RECT 31.530 107.985 31.760 108.220 ;
        RECT 33.110 107.985 33.340 108.220 ;
        RECT 35.150 107.985 35.380 108.230 ;
        RECT 36.730 107.985 36.960 108.230 ;
        RECT 38.040 108.220 38.770 112.570 ;
        RECT 39.620 108.220 40.350 112.570 ;
        RECT 41.210 108.220 41.940 112.570 ;
        RECT 42.780 108.220 43.510 112.570 ;
        RECT 43.750 111.390 44.500 111.450 ;
        RECT 43.730 108.970 44.520 111.390 ;
        RECT 43.750 108.910 44.500 108.970 ;
        RECT 44.690 108.230 45.420 112.580 ;
        RECT 46.280 108.230 47.010 112.580 ;
        RECT 48.110 112.570 48.340 117.985 ;
        RECT 49.690 112.570 49.920 117.985 ;
        RECT 51.270 112.570 51.500 117.985 ;
        RECT 52.850 112.570 53.080 117.985 ;
        RECT 38.310 107.985 38.540 108.220 ;
        RECT 39.890 107.985 40.120 108.220 ;
        RECT 41.470 107.985 41.700 108.220 ;
        RECT 43.050 107.985 43.280 108.220 ;
        RECT 44.950 107.985 45.180 108.230 ;
        RECT 46.530 107.985 46.760 108.230 ;
        RECT 47.850 108.220 48.580 112.570 ;
        RECT 49.430 108.220 50.160 112.570 ;
        RECT 51.020 108.220 51.750 112.570 ;
        RECT 52.590 108.220 53.320 112.570 ;
        RECT 54.750 112.550 54.980 117.985 ;
        RECT 56.330 112.550 56.560 117.985 ;
        RECT 48.110 107.985 48.340 108.220 ;
        RECT 49.690 107.985 49.920 108.220 ;
        RECT 51.270 107.985 51.500 108.220 ;
        RECT 52.850 107.985 53.080 108.220 ;
        RECT 54.500 108.200 55.230 112.550 ;
        RECT 56.090 108.200 56.820 112.550 ;
        RECT 57.910 112.540 58.140 117.985 ;
        RECT 59.490 112.540 59.720 117.985 ;
        RECT 61.070 112.540 61.300 117.985 ;
        RECT 62.650 112.540 62.880 117.985 ;
        RECT 64.550 112.550 64.780 117.985 ;
        RECT 66.130 112.550 66.360 117.985 ;
        RECT 54.750 107.985 54.980 108.200 ;
        RECT 56.330 107.985 56.560 108.200 ;
        RECT 57.660 108.190 58.390 112.540 ;
        RECT 59.240 108.190 59.970 112.540 ;
        RECT 60.830 108.190 61.560 112.540 ;
        RECT 62.400 108.190 63.130 112.540 ;
        RECT 63.330 111.370 64.080 111.430 ;
        RECT 63.310 108.950 64.100 111.370 ;
        RECT 63.330 108.890 64.080 108.950 ;
        RECT 64.290 108.200 65.020 112.550 ;
        RECT 65.880 108.200 66.610 112.550 ;
        RECT 67.710 112.540 67.940 117.985 ;
        RECT 69.290 112.540 69.520 117.985 ;
        RECT 70.870 112.540 71.100 117.985 ;
        RECT 72.450 112.540 72.680 117.985 ;
        RECT 57.910 107.985 58.140 108.190 ;
        RECT 59.490 107.985 59.720 108.190 ;
        RECT 61.070 107.985 61.300 108.190 ;
        RECT 62.650 107.985 62.880 108.190 ;
        RECT 64.550 107.985 64.780 108.200 ;
        RECT 66.130 107.985 66.360 108.200 ;
        RECT 67.450 108.190 68.180 112.540 ;
        RECT 69.030 108.190 69.760 112.540 ;
        RECT 70.620 108.190 71.350 112.540 ;
        RECT 72.190 108.190 72.920 112.540 ;
        RECT 67.710 107.985 67.940 108.190 ;
        RECT 69.290 107.985 69.520 108.190 ;
        RECT 70.870 107.985 71.100 108.190 ;
        RECT 72.450 107.985 72.680 108.190 ;
        RECT 25.210 101.400 25.440 106.805 ;
        RECT 26.790 101.400 27.020 106.805 ;
        RECT 24.950 97.050 25.680 101.400 ;
        RECT 26.540 97.050 27.270 101.400 ;
        RECT 28.370 101.390 28.600 106.805 ;
        RECT 29.950 101.390 30.180 106.805 ;
        RECT 31.530 101.390 31.760 106.805 ;
        RECT 33.110 101.390 33.340 106.805 ;
        RECT 35.150 101.400 35.380 106.805 ;
        RECT 36.730 101.400 36.960 106.805 ;
        RECT 25.210 96.805 25.440 97.050 ;
        RECT 26.790 96.805 27.020 97.050 ;
        RECT 28.110 97.040 28.840 101.390 ;
        RECT 29.690 97.040 30.420 101.390 ;
        RECT 31.280 97.040 32.010 101.390 ;
        RECT 32.850 97.040 33.580 101.390 ;
        RECT 33.840 100.450 34.590 100.510 ;
        RECT 33.820 98.030 34.610 100.450 ;
        RECT 33.840 97.970 34.590 98.030 ;
        RECT 34.880 97.050 35.610 101.400 ;
        RECT 36.470 97.050 37.200 101.400 ;
        RECT 38.310 101.390 38.540 106.805 ;
        RECT 39.890 101.390 40.120 106.805 ;
        RECT 41.470 101.390 41.700 106.805 ;
        RECT 43.050 101.390 43.280 106.805 ;
        RECT 44.950 101.400 45.180 106.805 ;
        RECT 46.530 101.400 46.760 106.805 ;
        RECT 28.370 96.805 28.600 97.040 ;
        RECT 29.950 96.805 30.180 97.040 ;
        RECT 31.530 96.805 31.760 97.040 ;
        RECT 33.110 96.805 33.340 97.040 ;
        RECT 35.150 96.805 35.380 97.050 ;
        RECT 36.730 96.805 36.960 97.050 ;
        RECT 38.040 97.040 38.770 101.390 ;
        RECT 39.620 97.040 40.350 101.390 ;
        RECT 41.210 97.040 41.940 101.390 ;
        RECT 42.780 97.040 43.510 101.390 ;
        RECT 44.690 97.050 45.420 101.400 ;
        RECT 46.280 97.050 47.010 101.400 ;
        RECT 48.110 101.390 48.340 106.805 ;
        RECT 49.690 101.390 49.920 106.805 ;
        RECT 51.270 101.390 51.500 106.805 ;
        RECT 52.850 101.390 53.080 106.805 ;
        RECT 38.310 96.805 38.540 97.040 ;
        RECT 39.890 96.805 40.120 97.040 ;
        RECT 41.470 96.805 41.700 97.040 ;
        RECT 43.050 96.805 43.280 97.040 ;
        RECT 44.950 96.805 45.180 97.050 ;
        RECT 46.530 96.805 46.760 97.050 ;
        RECT 47.850 97.040 48.580 101.390 ;
        RECT 49.430 97.040 50.160 101.390 ;
        RECT 51.020 97.040 51.750 101.390 ;
        RECT 52.590 97.040 53.320 101.390 ;
        RECT 54.750 101.370 54.980 106.805 ;
        RECT 56.330 101.370 56.560 106.805 ;
        RECT 53.570 100.410 54.320 100.470 ;
        RECT 53.550 97.990 54.340 100.410 ;
        RECT 53.570 97.930 54.320 97.990 ;
        RECT 48.110 96.805 48.340 97.040 ;
        RECT 49.690 96.805 49.920 97.040 ;
        RECT 51.270 96.805 51.500 97.040 ;
        RECT 52.850 96.805 53.080 97.040 ;
        RECT 54.500 97.020 55.230 101.370 ;
        RECT 56.090 97.020 56.820 101.370 ;
        RECT 57.910 101.360 58.140 106.805 ;
        RECT 59.490 101.360 59.720 106.805 ;
        RECT 61.070 101.360 61.300 106.805 ;
        RECT 62.650 101.360 62.880 106.805 ;
        RECT 64.550 101.370 64.780 106.805 ;
        RECT 66.130 101.370 66.360 106.805 ;
        RECT 54.750 96.805 54.980 97.020 ;
        RECT 56.330 96.805 56.560 97.020 ;
        RECT 57.660 97.010 58.390 101.360 ;
        RECT 59.240 97.010 59.970 101.360 ;
        RECT 60.830 97.010 61.560 101.360 ;
        RECT 62.400 97.010 63.130 101.360 ;
        RECT 64.290 97.020 65.020 101.370 ;
        RECT 65.880 97.020 66.610 101.370 ;
        RECT 67.710 101.360 67.940 106.805 ;
        RECT 69.290 101.360 69.520 106.805 ;
        RECT 70.870 101.360 71.100 106.805 ;
        RECT 72.450 101.360 72.680 106.805 ;
        RECT 57.910 96.805 58.140 97.010 ;
        RECT 59.490 96.805 59.720 97.010 ;
        RECT 61.070 96.805 61.300 97.010 ;
        RECT 62.650 96.805 62.880 97.010 ;
        RECT 64.550 96.805 64.780 97.020 ;
        RECT 66.130 96.805 66.360 97.020 ;
        RECT 67.450 97.010 68.180 101.360 ;
        RECT 69.030 97.010 69.760 101.360 ;
        RECT 70.620 97.010 71.350 101.360 ;
        RECT 72.190 97.010 72.920 101.360 ;
        RECT 67.710 96.805 67.940 97.010 ;
        RECT 69.290 96.805 69.520 97.010 ;
        RECT 70.870 96.805 71.100 97.010 ;
        RECT 72.450 96.805 72.680 97.010 ;
        RECT 7.905 80.455 8.235 80.515 ;
        RECT 3.255 79.855 3.645 80.455 ;
        RECT 4.835 79.855 5.225 80.455 ;
        RECT 6.415 79.855 6.805 80.455 ;
        RECT 7.885 79.855 8.255 80.455 ;
        RECT 9.335 79.855 9.725 80.455 ;
        RECT 10.915 79.855 11.305 80.455 ;
        RECT 12.495 79.855 12.885 80.455 ;
        RECT 3.335 78.450 3.565 79.855 ;
        RECT 4.915 78.450 5.145 79.855 ;
        RECT 6.495 78.450 6.725 79.855 ;
        RECT 7.905 79.795 8.235 79.855 ;
        RECT 9.415 78.450 9.645 79.855 ;
        RECT 10.995 78.450 11.225 79.855 ;
        RECT 12.575 78.450 12.805 79.855 ;
        RECT 17.705 79.800 17.935 79.870 ;
        RECT 19.285 79.800 19.515 79.870 ;
        RECT 19.915 79.800 20.395 79.860 ;
        RECT 20.785 79.800 21.015 79.870 ;
        RECT 22.365 79.800 22.595 79.870 ;
        RECT 17.645 78.950 18.005 79.800 ;
        RECT 19.225 78.950 19.585 79.800 ;
        RECT 19.895 78.950 20.415 79.800 ;
        RECT 20.725 78.950 21.085 79.800 ;
        RECT 22.305 78.950 22.665 79.800 ;
        RECT 17.705 69.870 17.935 78.950 ;
        RECT 19.285 69.870 19.515 78.950 ;
        RECT 19.915 78.890 20.395 78.950 ;
        RECT 20.785 69.870 21.015 78.950 ;
        RECT 22.365 69.870 22.595 78.950 ;
        RECT 1.270 28.260 1.500 56.485 ;
        RECT 11.560 28.260 11.790 56.485 ;
        RECT 25.210 44.780 25.440 45.025 ;
        RECT 26.790 44.780 27.020 45.025 ;
        RECT 28.370 44.790 28.600 45.025 ;
        RECT 29.950 44.790 30.180 45.025 ;
        RECT 31.530 44.790 31.760 45.025 ;
        RECT 33.110 44.790 33.340 45.025 ;
        RECT 24.950 40.430 25.680 44.780 ;
        RECT 26.540 40.430 27.270 44.780 ;
        RECT 28.110 40.440 28.840 44.790 ;
        RECT 29.690 40.440 30.420 44.790 ;
        RECT 31.280 40.440 32.010 44.790 ;
        RECT 32.850 40.440 33.580 44.790 ;
        RECT 35.150 44.780 35.380 45.025 ;
        RECT 36.730 44.780 36.960 45.025 ;
        RECT 38.310 44.790 38.540 45.025 ;
        RECT 39.890 44.790 40.120 45.025 ;
        RECT 41.470 44.790 41.700 45.025 ;
        RECT 43.050 44.790 43.280 45.025 ;
        RECT 33.840 43.800 34.590 43.860 ;
        RECT 33.820 41.380 34.610 43.800 ;
        RECT 33.840 41.320 34.590 41.380 ;
        RECT 17.065 32.610 17.295 32.810 ;
        RECT 16.980 31.960 17.380 32.610 ;
        RECT 17.065 31.810 17.295 31.960 ;
        RECT 1.250 18.400 11.830 28.260 ;
        RECT 16.280 26.520 16.510 29.250 ;
        RECT 17.860 26.520 18.090 29.250 ;
        RECT 16.200 25.870 16.600 26.520 ;
        RECT 17.760 25.870 18.160 26.520 ;
        RECT 19.765 26.480 19.995 35.245 ;
        RECT 21.345 26.510 21.575 35.245 ;
        RECT 22.925 26.510 23.155 35.245 ;
        RECT 25.210 35.025 25.440 40.430 ;
        RECT 26.790 35.025 27.020 40.430 ;
        RECT 28.370 35.025 28.600 40.440 ;
        RECT 29.950 35.025 30.180 40.440 ;
        RECT 31.530 35.025 31.760 40.440 ;
        RECT 33.110 35.025 33.340 40.440 ;
        RECT 34.880 40.430 35.610 44.780 ;
        RECT 36.470 40.430 37.200 44.780 ;
        RECT 38.040 40.440 38.770 44.790 ;
        RECT 39.620 40.440 40.350 44.790 ;
        RECT 41.210 40.440 41.940 44.790 ;
        RECT 42.780 40.440 43.510 44.790 ;
        RECT 44.950 44.780 45.180 45.025 ;
        RECT 46.530 44.780 46.760 45.025 ;
        RECT 48.110 44.790 48.340 45.025 ;
        RECT 49.690 44.790 49.920 45.025 ;
        RECT 51.270 44.790 51.500 45.025 ;
        RECT 52.850 44.790 53.080 45.025 ;
        RECT 54.750 44.810 54.980 45.025 ;
        RECT 56.330 44.810 56.560 45.025 ;
        RECT 57.910 44.820 58.140 45.025 ;
        RECT 59.490 44.820 59.720 45.025 ;
        RECT 61.070 44.820 61.300 45.025 ;
        RECT 62.650 44.820 62.880 45.025 ;
        RECT 35.150 35.025 35.380 40.430 ;
        RECT 36.730 35.025 36.960 40.430 ;
        RECT 38.310 35.025 38.540 40.440 ;
        RECT 39.890 35.025 40.120 40.440 ;
        RECT 41.470 35.025 41.700 40.440 ;
        RECT 43.050 35.025 43.280 40.440 ;
        RECT 44.690 40.430 45.420 44.780 ;
        RECT 46.280 40.430 47.010 44.780 ;
        RECT 47.850 40.440 48.580 44.790 ;
        RECT 49.430 40.440 50.160 44.790 ;
        RECT 51.020 40.440 51.750 44.790 ;
        RECT 52.590 40.440 53.320 44.790 ;
        RECT 53.570 43.840 54.320 43.900 ;
        RECT 53.550 41.420 54.340 43.840 ;
        RECT 53.570 41.360 54.320 41.420 ;
        RECT 54.500 40.460 55.230 44.810 ;
        RECT 56.090 40.460 56.820 44.810 ;
        RECT 57.660 40.470 58.390 44.820 ;
        RECT 59.240 40.470 59.970 44.820 ;
        RECT 60.830 40.470 61.560 44.820 ;
        RECT 62.400 40.470 63.130 44.820 ;
        RECT 64.550 44.810 64.780 45.025 ;
        RECT 66.130 44.810 66.360 45.025 ;
        RECT 67.710 44.820 67.940 45.025 ;
        RECT 69.290 44.820 69.520 45.025 ;
        RECT 70.870 44.820 71.100 45.025 ;
        RECT 72.450 44.820 72.680 45.025 ;
        RECT 44.950 35.025 45.180 40.430 ;
        RECT 46.530 35.025 46.760 40.430 ;
        RECT 48.110 35.025 48.340 40.440 ;
        RECT 49.690 35.025 49.920 40.440 ;
        RECT 51.270 35.025 51.500 40.440 ;
        RECT 52.850 35.025 53.080 40.440 ;
        RECT 54.750 35.025 54.980 40.460 ;
        RECT 56.330 35.025 56.560 40.460 ;
        RECT 57.910 35.025 58.140 40.470 ;
        RECT 59.490 35.025 59.720 40.470 ;
        RECT 61.070 35.025 61.300 40.470 ;
        RECT 62.650 35.025 62.880 40.470 ;
        RECT 64.290 40.460 65.020 44.810 ;
        RECT 65.880 40.460 66.610 44.810 ;
        RECT 67.450 40.470 68.180 44.820 ;
        RECT 69.030 40.470 69.760 44.820 ;
        RECT 70.620 40.470 71.350 44.820 ;
        RECT 72.190 40.470 72.920 44.820 ;
        RECT 64.550 35.025 64.780 40.460 ;
        RECT 66.130 35.025 66.360 40.460 ;
        RECT 67.710 35.025 67.940 40.470 ;
        RECT 69.290 35.025 69.520 40.470 ;
        RECT 70.870 35.025 71.100 40.470 ;
        RECT 72.450 35.025 72.680 40.470 ;
        RECT 25.210 33.600 25.440 33.845 ;
        RECT 26.790 33.600 27.020 33.845 ;
        RECT 28.370 33.610 28.600 33.845 ;
        RECT 29.950 33.610 30.180 33.845 ;
        RECT 31.530 33.610 31.760 33.845 ;
        RECT 33.110 33.610 33.340 33.845 ;
        RECT 24.950 29.250 25.680 33.600 ;
        RECT 26.540 29.250 27.270 33.600 ;
        RECT 28.110 29.260 28.840 33.610 ;
        RECT 29.690 29.260 30.420 33.610 ;
        RECT 31.280 29.260 32.010 33.610 ;
        RECT 32.850 29.260 33.580 33.610 ;
        RECT 35.150 33.600 35.380 33.845 ;
        RECT 36.730 33.600 36.960 33.845 ;
        RECT 38.310 33.610 38.540 33.845 ;
        RECT 39.890 33.610 40.120 33.845 ;
        RECT 41.470 33.610 41.700 33.845 ;
        RECT 43.050 33.610 43.280 33.845 ;
        RECT 16.280 25.250 16.510 25.870 ;
        RECT 17.860 25.250 18.090 25.870 ;
        RECT 19.670 25.830 20.070 26.480 ;
        RECT 21.260 25.860 21.660 26.510 ;
        RECT 22.820 25.860 23.220 26.510 ;
        RECT 19.765 25.245 19.995 25.830 ;
        RECT 21.345 25.245 21.575 25.860 ;
        RECT 22.925 25.245 23.155 25.860 ;
        RECT 25.210 23.845 25.440 29.250 ;
        RECT 26.790 23.845 27.020 29.250 ;
        RECT 28.370 23.845 28.600 29.260 ;
        RECT 29.950 23.845 30.180 29.260 ;
        RECT 31.530 23.845 31.760 29.260 ;
        RECT 33.110 23.845 33.340 29.260 ;
        RECT 34.880 29.250 35.610 33.600 ;
        RECT 36.470 29.250 37.200 33.600 ;
        RECT 38.040 29.260 38.770 33.610 ;
        RECT 39.620 29.260 40.350 33.610 ;
        RECT 41.210 29.260 41.940 33.610 ;
        RECT 42.780 29.260 43.510 33.610 ;
        RECT 44.950 33.600 45.180 33.845 ;
        RECT 46.530 33.600 46.760 33.845 ;
        RECT 48.110 33.610 48.340 33.845 ;
        RECT 49.690 33.610 49.920 33.845 ;
        RECT 51.270 33.610 51.500 33.845 ;
        RECT 52.850 33.610 53.080 33.845 ;
        RECT 54.750 33.630 54.980 33.845 ;
        RECT 56.330 33.630 56.560 33.845 ;
        RECT 57.910 33.640 58.140 33.845 ;
        RECT 59.490 33.640 59.720 33.845 ;
        RECT 61.070 33.640 61.300 33.845 ;
        RECT 62.650 33.640 62.880 33.845 ;
        RECT 43.750 32.860 44.500 32.920 ;
        RECT 43.730 30.440 44.520 32.860 ;
        RECT 43.750 30.380 44.500 30.440 ;
        RECT 35.150 23.845 35.380 29.250 ;
        RECT 36.730 23.845 36.960 29.250 ;
        RECT 38.310 23.845 38.540 29.260 ;
        RECT 39.890 23.845 40.120 29.260 ;
        RECT 41.470 23.845 41.700 29.260 ;
        RECT 43.050 23.845 43.280 29.260 ;
        RECT 44.690 29.250 45.420 33.600 ;
        RECT 46.280 29.250 47.010 33.600 ;
        RECT 47.850 29.260 48.580 33.610 ;
        RECT 49.430 29.260 50.160 33.610 ;
        RECT 51.020 29.260 51.750 33.610 ;
        RECT 52.590 29.260 53.320 33.610 ;
        RECT 54.500 29.280 55.230 33.630 ;
        RECT 56.090 29.280 56.820 33.630 ;
        RECT 57.660 29.290 58.390 33.640 ;
        RECT 59.240 29.290 59.970 33.640 ;
        RECT 60.830 29.290 61.560 33.640 ;
        RECT 62.400 29.290 63.130 33.640 ;
        RECT 64.550 33.630 64.780 33.845 ;
        RECT 66.130 33.630 66.360 33.845 ;
        RECT 67.710 33.640 67.940 33.845 ;
        RECT 69.290 33.640 69.520 33.845 ;
        RECT 70.870 33.640 71.100 33.845 ;
        RECT 72.450 33.640 72.680 33.845 ;
        RECT 63.330 32.880 64.080 32.940 ;
        RECT 63.310 30.460 64.100 32.880 ;
        RECT 63.330 30.400 64.080 30.460 ;
        RECT 44.950 23.845 45.180 29.250 ;
        RECT 46.530 23.845 46.760 29.250 ;
        RECT 48.110 23.845 48.340 29.260 ;
        RECT 49.690 23.845 49.920 29.260 ;
        RECT 51.270 23.845 51.500 29.260 ;
        RECT 52.850 23.845 53.080 29.260 ;
        RECT 54.750 23.845 54.980 29.280 ;
        RECT 56.330 23.845 56.560 29.280 ;
        RECT 57.910 23.845 58.140 29.290 ;
        RECT 59.490 23.845 59.720 29.290 ;
        RECT 61.070 23.845 61.300 29.290 ;
        RECT 62.650 23.845 62.880 29.290 ;
        RECT 64.290 29.280 65.020 33.630 ;
        RECT 65.880 29.280 66.610 33.630 ;
        RECT 67.450 29.290 68.180 33.640 ;
        RECT 69.030 29.290 69.760 33.640 ;
        RECT 70.620 29.290 71.350 33.640 ;
        RECT 72.190 29.290 72.920 33.640 ;
        RECT 64.550 23.845 64.780 29.280 ;
        RECT 66.130 23.845 66.360 29.280 ;
        RECT 67.710 23.845 67.940 29.290 ;
        RECT 69.290 23.845 69.520 29.290 ;
        RECT 70.870 23.845 71.100 29.290 ;
        RECT 72.450 23.845 72.680 29.290 ;
        RECT 15.025 22.010 15.255 22.665 ;
        RECT 14.930 21.360 15.330 22.010 ;
        RECT 16.605 22.000 16.835 22.665 ;
        RECT 18.185 22.010 18.415 22.665 ;
        RECT 19.765 22.020 19.995 22.665 ;
        RECT 21.345 22.020 21.575 22.665 ;
        RECT 22.925 22.020 23.155 22.665 ;
        RECT 25.210 22.420 25.440 22.665 ;
        RECT 26.790 22.420 27.020 22.665 ;
        RECT 28.370 22.430 28.600 22.665 ;
        RECT 29.950 22.430 30.180 22.665 ;
        RECT 31.530 22.430 31.760 22.665 ;
        RECT 33.110 22.430 33.340 22.665 ;
        RECT 1.270 1.485 1.500 18.400 ;
        RECT 11.560 1.485 11.790 18.400 ;
        RECT 15.025 12.665 15.255 21.360 ;
        RECT 16.510 21.350 16.910 22.000 ;
        RECT 18.080 21.360 18.480 22.010 ;
        RECT 19.680 21.370 20.080 22.020 ;
        RECT 21.260 21.370 21.660 22.020 ;
        RECT 22.840 21.370 23.240 22.020 ;
        RECT 16.605 12.665 16.835 21.350 ;
        RECT 18.185 12.665 18.415 21.360 ;
        RECT 19.765 12.665 19.995 21.370 ;
        RECT 21.345 12.665 21.575 21.370 ;
        RECT 22.925 12.665 23.155 21.370 ;
        RECT 24.950 18.070 25.680 22.420 ;
        RECT 26.540 18.070 27.270 22.420 ;
        RECT 28.110 18.080 28.840 22.430 ;
        RECT 29.690 18.080 30.420 22.430 ;
        RECT 31.280 18.080 32.010 22.430 ;
        RECT 32.850 18.080 33.580 22.430 ;
        RECT 35.150 22.420 35.380 22.665 ;
        RECT 36.730 22.420 36.960 22.665 ;
        RECT 38.310 22.430 38.540 22.665 ;
        RECT 39.890 22.430 40.120 22.665 ;
        RECT 41.470 22.430 41.700 22.665 ;
        RECT 43.050 22.430 43.280 22.665 ;
        RECT 33.860 21.610 34.610 21.670 ;
        RECT 33.840 19.190 34.630 21.610 ;
        RECT 33.860 19.130 34.610 19.190 ;
        RECT 25.210 12.665 25.440 18.070 ;
        RECT 26.790 12.665 27.020 18.070 ;
        RECT 28.370 12.665 28.600 18.080 ;
        RECT 29.950 12.665 30.180 18.080 ;
        RECT 31.530 12.665 31.760 18.080 ;
        RECT 33.110 12.665 33.340 18.080 ;
        RECT 34.880 18.070 35.610 22.420 ;
        RECT 36.470 18.070 37.200 22.420 ;
        RECT 38.040 18.080 38.770 22.430 ;
        RECT 39.620 18.080 40.350 22.430 ;
        RECT 41.210 18.080 41.940 22.430 ;
        RECT 42.780 18.080 43.510 22.430 ;
        RECT 44.950 22.420 45.180 22.665 ;
        RECT 46.530 22.420 46.760 22.665 ;
        RECT 48.110 22.430 48.340 22.665 ;
        RECT 49.690 22.430 49.920 22.665 ;
        RECT 51.270 22.430 51.500 22.665 ;
        RECT 52.850 22.430 53.080 22.665 ;
        RECT 54.750 22.450 54.980 22.665 ;
        RECT 56.330 22.450 56.560 22.665 ;
        RECT 57.910 22.460 58.140 22.665 ;
        RECT 59.490 22.460 59.720 22.665 ;
        RECT 61.070 22.460 61.300 22.665 ;
        RECT 62.650 22.460 62.880 22.665 ;
        RECT 35.150 12.665 35.380 18.070 ;
        RECT 36.730 12.665 36.960 18.070 ;
        RECT 38.310 12.665 38.540 18.080 ;
        RECT 39.890 12.665 40.120 18.080 ;
        RECT 41.470 12.665 41.700 18.080 ;
        RECT 43.050 12.665 43.280 18.080 ;
        RECT 44.690 18.070 45.420 22.420 ;
        RECT 46.280 18.070 47.010 22.420 ;
        RECT 47.850 18.080 48.580 22.430 ;
        RECT 49.430 18.080 50.160 22.430 ;
        RECT 51.020 18.080 51.750 22.430 ;
        RECT 52.590 18.080 53.320 22.430 ;
        RECT 53.540 21.610 54.290 21.670 ;
        RECT 53.520 19.190 54.310 21.610 ;
        RECT 53.540 19.130 54.290 19.190 ;
        RECT 54.500 18.100 55.230 22.450 ;
        RECT 56.090 18.100 56.820 22.450 ;
        RECT 57.660 18.110 58.390 22.460 ;
        RECT 59.240 18.110 59.970 22.460 ;
        RECT 60.830 18.110 61.560 22.460 ;
        RECT 62.400 18.110 63.130 22.460 ;
        RECT 64.550 22.450 64.780 22.665 ;
        RECT 66.130 22.450 66.360 22.665 ;
        RECT 67.710 22.460 67.940 22.665 ;
        RECT 69.290 22.460 69.520 22.665 ;
        RECT 70.870 22.460 71.100 22.665 ;
        RECT 72.450 22.460 72.680 22.665 ;
        RECT 44.950 12.665 45.180 18.070 ;
        RECT 46.530 12.665 46.760 18.070 ;
        RECT 48.110 12.665 48.340 18.080 ;
        RECT 49.690 12.665 49.920 18.080 ;
        RECT 51.270 12.665 51.500 18.080 ;
        RECT 52.850 12.665 53.080 18.080 ;
        RECT 54.750 12.665 54.980 18.100 ;
        RECT 56.330 12.665 56.560 18.100 ;
        RECT 57.910 12.665 58.140 18.110 ;
        RECT 59.490 12.665 59.720 18.110 ;
        RECT 61.070 12.665 61.300 18.110 ;
        RECT 62.650 12.665 62.880 18.110 ;
        RECT 64.290 18.100 65.020 22.450 ;
        RECT 65.880 18.100 66.610 22.450 ;
        RECT 67.450 18.110 68.180 22.460 ;
        RECT 69.030 18.110 69.760 22.460 ;
        RECT 70.620 18.110 71.350 22.460 ;
        RECT 72.190 18.110 72.920 22.460 ;
        RECT 64.550 12.665 64.780 18.100 ;
        RECT 66.130 12.665 66.360 18.100 ;
        RECT 67.710 12.665 67.940 18.110 ;
        RECT 69.290 12.665 69.520 18.110 ;
        RECT 70.870 12.665 71.100 18.110 ;
        RECT 72.450 12.665 72.680 18.110 ;
        RECT 15.025 2.610 15.255 11.485 ;
        RECT 14.950 1.960 15.350 2.610 ;
        RECT 16.605 2.600 16.835 11.485 ;
        RECT 18.185 2.610 18.415 11.485 ;
        RECT 15.025 1.485 15.255 1.960 ;
        RECT 16.510 1.950 16.910 2.600 ;
        RECT 18.110 1.960 18.510 2.610 ;
        RECT 19.765 2.600 19.995 11.485 ;
        RECT 21.345 2.610 21.575 11.485 ;
        RECT 22.925 2.610 23.155 11.485 ;
        RECT 25.210 11.240 25.440 11.485 ;
        RECT 26.790 11.240 27.020 11.485 ;
        RECT 28.370 11.250 28.600 11.485 ;
        RECT 29.950 11.250 30.180 11.485 ;
        RECT 31.530 11.250 31.760 11.485 ;
        RECT 33.110 11.250 33.340 11.485 ;
        RECT 24.950 6.890 25.680 11.240 ;
        RECT 26.540 6.890 27.270 11.240 ;
        RECT 28.110 6.900 28.840 11.250 ;
        RECT 29.690 6.900 30.420 11.250 ;
        RECT 31.280 6.900 32.010 11.250 ;
        RECT 32.850 6.900 33.580 11.250 ;
        RECT 35.150 11.240 35.380 11.485 ;
        RECT 36.730 11.240 36.960 11.485 ;
        RECT 38.310 11.250 38.540 11.485 ;
        RECT 39.890 11.250 40.120 11.485 ;
        RECT 41.470 11.250 41.700 11.485 ;
        RECT 43.050 11.250 43.280 11.485 ;
        RECT 16.605 1.485 16.835 1.950 ;
        RECT 18.185 1.485 18.415 1.960 ;
        RECT 19.680 1.950 20.080 2.600 ;
        RECT 21.260 1.960 21.660 2.610 ;
        RECT 22.840 1.960 23.240 2.610 ;
        RECT 19.765 1.485 19.995 1.950 ;
        RECT 21.345 1.485 21.575 1.960 ;
        RECT 22.925 1.485 23.155 1.960 ;
        RECT 25.210 1.485 25.440 6.890 ;
        RECT 26.790 1.485 27.020 6.890 ;
        RECT 28.370 1.485 28.600 6.900 ;
        RECT 29.950 1.485 30.180 6.900 ;
        RECT 31.530 1.485 31.760 6.900 ;
        RECT 33.110 1.485 33.340 6.900 ;
        RECT 34.880 6.890 35.610 11.240 ;
        RECT 36.470 6.890 37.200 11.240 ;
        RECT 38.040 6.900 38.770 11.250 ;
        RECT 39.620 6.900 40.350 11.250 ;
        RECT 41.210 6.900 41.940 11.250 ;
        RECT 42.780 6.900 43.510 11.250 ;
        RECT 44.950 11.240 45.180 11.485 ;
        RECT 46.530 11.240 46.760 11.485 ;
        RECT 48.110 11.250 48.340 11.485 ;
        RECT 49.690 11.250 49.920 11.485 ;
        RECT 51.270 11.250 51.500 11.485 ;
        RECT 52.850 11.250 53.080 11.485 ;
        RECT 54.750 11.270 54.980 11.485 ;
        RECT 56.330 11.270 56.560 11.485 ;
        RECT 57.910 11.280 58.140 11.485 ;
        RECT 59.490 11.280 59.720 11.485 ;
        RECT 61.070 11.280 61.300 11.485 ;
        RECT 62.650 11.280 62.880 11.485 ;
        RECT 43.760 10.470 44.510 10.530 ;
        RECT 43.740 8.050 44.530 10.470 ;
        RECT 43.760 7.990 44.510 8.050 ;
        RECT 35.150 1.485 35.380 6.890 ;
        RECT 36.730 1.485 36.960 6.890 ;
        RECT 38.310 1.485 38.540 6.900 ;
        RECT 39.890 1.485 40.120 6.900 ;
        RECT 41.470 1.485 41.700 6.900 ;
        RECT 43.050 1.485 43.280 6.900 ;
        RECT 44.690 6.890 45.420 11.240 ;
        RECT 46.280 6.890 47.010 11.240 ;
        RECT 47.850 6.900 48.580 11.250 ;
        RECT 49.430 6.900 50.160 11.250 ;
        RECT 51.020 6.900 51.750 11.250 ;
        RECT 52.590 6.900 53.320 11.250 ;
        RECT 54.500 6.920 55.230 11.270 ;
        RECT 56.090 6.920 56.820 11.270 ;
        RECT 57.660 6.930 58.390 11.280 ;
        RECT 59.240 6.930 59.970 11.280 ;
        RECT 60.830 6.930 61.560 11.280 ;
        RECT 62.400 6.930 63.130 11.280 ;
        RECT 64.550 11.270 64.780 11.485 ;
        RECT 66.130 11.270 66.360 11.485 ;
        RECT 67.710 11.280 67.940 11.485 ;
        RECT 69.290 11.280 69.520 11.485 ;
        RECT 70.870 11.280 71.100 11.485 ;
        RECT 72.450 11.280 72.680 11.485 ;
        RECT 63.320 10.430 64.070 10.490 ;
        RECT 63.300 8.010 64.090 10.430 ;
        RECT 63.320 7.950 64.070 8.010 ;
        RECT 44.950 1.485 45.180 6.890 ;
        RECT 46.530 1.485 46.760 6.890 ;
        RECT 48.110 1.485 48.340 6.900 ;
        RECT 49.690 1.485 49.920 6.900 ;
        RECT 51.270 1.485 51.500 6.900 ;
        RECT 52.850 1.485 53.080 6.900 ;
        RECT 54.750 1.485 54.980 6.920 ;
        RECT 56.330 1.485 56.560 6.920 ;
        RECT 57.910 1.485 58.140 6.930 ;
        RECT 59.490 1.485 59.720 6.930 ;
        RECT 61.070 1.485 61.300 6.930 ;
        RECT 62.650 1.485 62.880 6.930 ;
        RECT 64.290 6.920 65.020 11.270 ;
        RECT 65.880 6.920 66.610 11.270 ;
        RECT 67.450 6.930 68.180 11.280 ;
        RECT 69.030 6.930 69.760 11.280 ;
        RECT 70.620 6.930 71.350 11.280 ;
        RECT 72.190 6.930 72.920 11.280 ;
        RECT 64.550 1.485 64.780 6.920 ;
        RECT 66.130 1.485 66.360 6.920 ;
        RECT 67.710 1.485 67.940 6.930 ;
        RECT 69.290 1.485 69.520 6.930 ;
        RECT 70.870 1.485 71.100 6.930 ;
        RECT 72.450 1.485 72.680 6.930 ;
      LAYER via ;
        RECT 15.000 139.220 15.300 139.870 ;
        RECT 16.560 139.230 16.860 139.880 ;
        RECT 18.160 139.220 18.460 139.870 ;
        RECT 19.730 139.230 20.030 139.880 ;
        RECT 21.310 139.220 21.610 139.870 ;
        RECT 22.890 139.220 23.190 139.870 ;
        RECT 25.000 130.590 25.630 134.940 ;
        RECT 26.590 130.590 27.220 134.940 ;
        RECT 28.160 130.580 28.790 134.930 ;
        RECT 29.740 130.580 30.370 134.930 ;
        RECT 31.330 130.580 31.960 134.930 ;
        RECT 32.900 130.580 33.530 134.930 ;
        RECT 34.930 130.590 35.560 134.940 ;
        RECT 36.520 130.590 37.150 134.940 ;
        RECT 38.090 130.580 38.720 134.930 ;
        RECT 39.670 130.580 40.300 134.930 ;
        RECT 41.260 130.580 41.890 134.930 ;
        RECT 42.830 130.580 43.460 134.930 ;
        RECT 43.790 131.360 44.480 133.780 ;
        RECT 44.740 130.590 45.370 134.940 ;
        RECT 46.330 130.590 46.960 134.940 ;
        RECT 47.900 130.580 48.530 134.930 ;
        RECT 49.480 130.580 50.110 134.930 ;
        RECT 51.070 130.580 51.700 134.930 ;
        RECT 52.640 130.580 53.270 134.930 ;
        RECT 54.550 130.560 55.180 134.910 ;
        RECT 56.140 130.560 56.770 134.910 ;
        RECT 57.710 130.550 58.340 134.900 ;
        RECT 59.290 130.550 59.920 134.900 ;
        RECT 60.880 130.550 61.510 134.900 ;
        RECT 62.450 130.550 63.080 134.900 ;
        RECT 63.350 131.400 64.040 133.820 ;
        RECT 64.340 130.560 64.970 134.910 ;
        RECT 65.930 130.560 66.560 134.910 ;
        RECT 67.500 130.550 68.130 134.900 ;
        RECT 69.080 130.550 69.710 134.900 ;
        RECT 70.670 130.550 71.300 134.900 ;
        RECT 72.240 130.550 72.870 134.900 ;
        RECT 1.440 116.030 11.810 126.160 ;
        RECT 14.980 119.820 15.280 120.470 ;
        RECT 16.560 119.830 16.860 120.480 ;
        RECT 18.130 119.820 18.430 120.470 ;
        RECT 19.730 119.810 20.030 120.460 ;
        RECT 21.310 119.810 21.610 120.460 ;
        RECT 22.890 119.810 23.190 120.460 ;
        RECT 25.000 119.410 25.630 123.760 ;
        RECT 26.590 119.410 27.220 123.760 ;
        RECT 28.160 119.400 28.790 123.750 ;
        RECT 29.740 119.400 30.370 123.750 ;
        RECT 31.330 119.400 31.960 123.750 ;
        RECT 32.900 119.400 33.530 123.750 ;
        RECT 33.890 120.220 34.580 122.640 ;
        RECT 34.930 119.410 35.560 123.760 ;
        RECT 36.520 119.410 37.150 123.760 ;
        RECT 38.090 119.400 38.720 123.750 ;
        RECT 39.670 119.400 40.300 123.750 ;
        RECT 41.260 119.400 41.890 123.750 ;
        RECT 42.830 119.400 43.460 123.750 ;
        RECT 44.740 119.410 45.370 123.760 ;
        RECT 46.330 119.410 46.960 123.760 ;
        RECT 47.900 119.400 48.530 123.750 ;
        RECT 49.480 119.400 50.110 123.750 ;
        RECT 51.070 119.400 51.700 123.750 ;
        RECT 52.640 119.400 53.270 123.750 ;
        RECT 53.570 120.220 54.260 122.640 ;
        RECT 54.550 119.380 55.180 123.730 ;
        RECT 56.140 119.380 56.770 123.730 ;
        RECT 57.710 119.370 58.340 123.720 ;
        RECT 59.290 119.370 59.920 123.720 ;
        RECT 60.880 119.370 61.510 123.720 ;
        RECT 62.450 119.370 63.080 123.720 ;
        RECT 64.340 119.380 64.970 123.730 ;
        RECT 65.930 119.380 66.560 123.730 ;
        RECT 67.500 119.370 68.130 123.720 ;
        RECT 69.080 119.370 69.710 123.720 ;
        RECT 70.670 119.370 71.300 123.720 ;
        RECT 72.240 119.370 72.870 123.720 ;
        RECT 16.250 115.310 16.550 115.960 ;
        RECT 17.810 115.310 18.110 115.960 ;
        RECT 19.720 115.350 20.020 116.000 ;
        RECT 17.030 109.220 17.330 109.870 ;
        RECT 21.310 115.320 21.610 115.970 ;
        RECT 22.870 115.320 23.170 115.970 ;
        RECT 25.000 108.230 25.630 112.580 ;
        RECT 26.590 108.230 27.220 112.580 ;
        RECT 28.160 108.220 28.790 112.570 ;
        RECT 29.740 108.220 30.370 112.570 ;
        RECT 31.330 108.220 31.960 112.570 ;
        RECT 32.900 108.220 33.530 112.570 ;
        RECT 34.930 108.230 35.560 112.580 ;
        RECT 36.520 108.230 37.150 112.580 ;
        RECT 38.090 108.220 38.720 112.570 ;
        RECT 39.670 108.220 40.300 112.570 ;
        RECT 41.260 108.220 41.890 112.570 ;
        RECT 42.830 108.220 43.460 112.570 ;
        RECT 43.780 108.970 44.470 111.390 ;
        RECT 44.740 108.230 45.370 112.580 ;
        RECT 46.330 108.230 46.960 112.580 ;
        RECT 47.900 108.220 48.530 112.570 ;
        RECT 49.480 108.220 50.110 112.570 ;
        RECT 51.070 108.220 51.700 112.570 ;
        RECT 52.640 108.220 53.270 112.570 ;
        RECT 54.550 108.200 55.180 112.550 ;
        RECT 56.140 108.200 56.770 112.550 ;
        RECT 57.710 108.190 58.340 112.540 ;
        RECT 59.290 108.190 59.920 112.540 ;
        RECT 60.880 108.190 61.510 112.540 ;
        RECT 62.450 108.190 63.080 112.540 ;
        RECT 63.360 108.950 64.050 111.370 ;
        RECT 64.340 108.200 64.970 112.550 ;
        RECT 65.930 108.200 66.560 112.550 ;
        RECT 67.500 108.190 68.130 112.540 ;
        RECT 69.080 108.190 69.710 112.540 ;
        RECT 70.670 108.190 71.300 112.540 ;
        RECT 72.240 108.190 72.870 112.540 ;
        RECT 25.000 97.050 25.630 101.400 ;
        RECT 26.590 97.050 27.220 101.400 ;
        RECT 28.160 97.040 28.790 101.390 ;
        RECT 29.740 97.040 30.370 101.390 ;
        RECT 31.330 97.040 31.960 101.390 ;
        RECT 32.900 97.040 33.530 101.390 ;
        RECT 33.870 98.030 34.560 100.450 ;
        RECT 34.930 97.050 35.560 101.400 ;
        RECT 36.520 97.050 37.150 101.400 ;
        RECT 38.090 97.040 38.720 101.390 ;
        RECT 39.670 97.040 40.300 101.390 ;
        RECT 41.260 97.040 41.890 101.390 ;
        RECT 42.830 97.040 43.460 101.390 ;
        RECT 44.740 97.050 45.370 101.400 ;
        RECT 46.330 97.050 46.960 101.400 ;
        RECT 47.900 97.040 48.530 101.390 ;
        RECT 49.480 97.040 50.110 101.390 ;
        RECT 51.070 97.040 51.700 101.390 ;
        RECT 52.640 97.040 53.270 101.390 ;
        RECT 53.600 97.990 54.290 100.410 ;
        RECT 54.550 97.020 55.180 101.370 ;
        RECT 56.140 97.020 56.770 101.370 ;
        RECT 57.710 97.010 58.340 101.360 ;
        RECT 59.290 97.010 59.920 101.360 ;
        RECT 60.880 97.010 61.510 101.360 ;
        RECT 62.450 97.010 63.080 101.360 ;
        RECT 64.340 97.020 64.970 101.370 ;
        RECT 65.930 97.020 66.560 101.370 ;
        RECT 67.500 97.010 68.130 101.360 ;
        RECT 69.080 97.010 69.710 101.360 ;
        RECT 70.670 97.010 71.300 101.360 ;
        RECT 72.240 97.010 72.870 101.360 ;
        RECT 3.305 79.855 3.595 80.455 ;
        RECT 4.885 79.855 5.175 80.455 ;
        RECT 6.465 79.855 6.755 80.455 ;
        RECT 7.935 79.855 8.205 80.455 ;
        RECT 9.385 79.855 9.675 80.455 ;
        RECT 10.965 79.855 11.255 80.455 ;
        RECT 12.545 79.855 12.835 80.455 ;
        RECT 17.695 78.950 17.955 79.800 ;
        RECT 19.275 78.950 19.535 79.800 ;
        RECT 19.945 78.950 20.365 79.800 ;
        RECT 20.775 78.950 21.035 79.800 ;
        RECT 22.355 78.950 22.615 79.800 ;
        RECT 25.000 40.430 25.630 44.780 ;
        RECT 26.590 40.430 27.220 44.780 ;
        RECT 28.160 40.440 28.790 44.790 ;
        RECT 29.740 40.440 30.370 44.790 ;
        RECT 31.330 40.440 31.960 44.790 ;
        RECT 32.900 40.440 33.530 44.790 ;
        RECT 33.870 41.380 34.560 43.800 ;
        RECT 17.030 31.960 17.330 32.610 ;
        RECT 1.300 18.400 11.780 28.260 ;
        RECT 16.250 25.870 16.550 26.520 ;
        RECT 17.810 25.870 18.110 26.520 ;
        RECT 34.930 40.430 35.560 44.780 ;
        RECT 36.520 40.430 37.150 44.780 ;
        RECT 38.090 40.440 38.720 44.790 ;
        RECT 39.670 40.440 40.300 44.790 ;
        RECT 41.260 40.440 41.890 44.790 ;
        RECT 42.830 40.440 43.460 44.790 ;
        RECT 44.740 40.430 45.370 44.780 ;
        RECT 46.330 40.430 46.960 44.780 ;
        RECT 47.900 40.440 48.530 44.790 ;
        RECT 49.480 40.440 50.110 44.790 ;
        RECT 51.070 40.440 51.700 44.790 ;
        RECT 52.640 40.440 53.270 44.790 ;
        RECT 53.600 41.420 54.290 43.840 ;
        RECT 54.550 40.460 55.180 44.810 ;
        RECT 56.140 40.460 56.770 44.810 ;
        RECT 57.710 40.470 58.340 44.820 ;
        RECT 59.290 40.470 59.920 44.820 ;
        RECT 60.880 40.470 61.510 44.820 ;
        RECT 62.450 40.470 63.080 44.820 ;
        RECT 64.340 40.460 64.970 44.810 ;
        RECT 65.930 40.460 66.560 44.810 ;
        RECT 67.500 40.470 68.130 44.820 ;
        RECT 69.080 40.470 69.710 44.820 ;
        RECT 70.670 40.470 71.300 44.820 ;
        RECT 72.240 40.470 72.870 44.820 ;
        RECT 25.000 29.250 25.630 33.600 ;
        RECT 26.590 29.250 27.220 33.600 ;
        RECT 28.160 29.260 28.790 33.610 ;
        RECT 29.740 29.260 30.370 33.610 ;
        RECT 31.330 29.260 31.960 33.610 ;
        RECT 32.900 29.260 33.530 33.610 ;
        RECT 19.720 25.830 20.020 26.480 ;
        RECT 21.310 25.860 21.610 26.510 ;
        RECT 22.870 25.860 23.170 26.510 ;
        RECT 34.930 29.250 35.560 33.600 ;
        RECT 36.520 29.250 37.150 33.600 ;
        RECT 38.090 29.260 38.720 33.610 ;
        RECT 39.670 29.260 40.300 33.610 ;
        RECT 41.260 29.260 41.890 33.610 ;
        RECT 42.830 29.260 43.460 33.610 ;
        RECT 43.780 30.440 44.470 32.860 ;
        RECT 44.740 29.250 45.370 33.600 ;
        RECT 46.330 29.250 46.960 33.600 ;
        RECT 47.900 29.260 48.530 33.610 ;
        RECT 49.480 29.260 50.110 33.610 ;
        RECT 51.070 29.260 51.700 33.610 ;
        RECT 52.640 29.260 53.270 33.610 ;
        RECT 54.550 29.280 55.180 33.630 ;
        RECT 56.140 29.280 56.770 33.630 ;
        RECT 57.710 29.290 58.340 33.640 ;
        RECT 59.290 29.290 59.920 33.640 ;
        RECT 60.880 29.290 61.510 33.640 ;
        RECT 62.450 29.290 63.080 33.640 ;
        RECT 63.360 30.460 64.050 32.880 ;
        RECT 64.340 29.280 64.970 33.630 ;
        RECT 65.930 29.280 66.560 33.630 ;
        RECT 67.500 29.290 68.130 33.640 ;
        RECT 69.080 29.290 69.710 33.640 ;
        RECT 70.670 29.290 71.300 33.640 ;
        RECT 72.240 29.290 72.870 33.640 ;
        RECT 14.980 21.360 15.280 22.010 ;
        RECT 16.560 21.350 16.860 22.000 ;
        RECT 18.130 21.360 18.430 22.010 ;
        RECT 19.730 21.370 20.030 22.020 ;
        RECT 21.310 21.370 21.610 22.020 ;
        RECT 22.890 21.370 23.190 22.020 ;
        RECT 25.000 18.070 25.630 22.420 ;
        RECT 26.590 18.070 27.220 22.420 ;
        RECT 28.160 18.080 28.790 22.430 ;
        RECT 29.740 18.080 30.370 22.430 ;
        RECT 31.330 18.080 31.960 22.430 ;
        RECT 32.900 18.080 33.530 22.430 ;
        RECT 33.890 19.190 34.580 21.610 ;
        RECT 34.930 18.070 35.560 22.420 ;
        RECT 36.520 18.070 37.150 22.420 ;
        RECT 38.090 18.080 38.720 22.430 ;
        RECT 39.670 18.080 40.300 22.430 ;
        RECT 41.260 18.080 41.890 22.430 ;
        RECT 42.830 18.080 43.460 22.430 ;
        RECT 44.740 18.070 45.370 22.420 ;
        RECT 46.330 18.070 46.960 22.420 ;
        RECT 47.900 18.080 48.530 22.430 ;
        RECT 49.480 18.080 50.110 22.430 ;
        RECT 51.070 18.080 51.700 22.430 ;
        RECT 52.640 18.080 53.270 22.430 ;
        RECT 53.570 19.190 54.260 21.610 ;
        RECT 54.550 18.100 55.180 22.450 ;
        RECT 56.140 18.100 56.770 22.450 ;
        RECT 57.710 18.110 58.340 22.460 ;
        RECT 59.290 18.110 59.920 22.460 ;
        RECT 60.880 18.110 61.510 22.460 ;
        RECT 62.450 18.110 63.080 22.460 ;
        RECT 64.340 18.100 64.970 22.450 ;
        RECT 65.930 18.100 66.560 22.450 ;
        RECT 67.500 18.110 68.130 22.460 ;
        RECT 69.080 18.110 69.710 22.460 ;
        RECT 70.670 18.110 71.300 22.460 ;
        RECT 72.240 18.110 72.870 22.460 ;
        RECT 15.000 1.960 15.300 2.610 ;
        RECT 16.560 1.950 16.860 2.600 ;
        RECT 18.160 1.960 18.460 2.610 ;
        RECT 25.000 6.890 25.630 11.240 ;
        RECT 26.590 6.890 27.220 11.240 ;
        RECT 28.160 6.900 28.790 11.250 ;
        RECT 29.740 6.900 30.370 11.250 ;
        RECT 31.330 6.900 31.960 11.250 ;
        RECT 32.900 6.900 33.530 11.250 ;
        RECT 19.730 1.950 20.030 2.600 ;
        RECT 21.310 1.960 21.610 2.610 ;
        RECT 22.890 1.960 23.190 2.610 ;
        RECT 34.930 6.890 35.560 11.240 ;
        RECT 36.520 6.890 37.150 11.240 ;
        RECT 38.090 6.900 38.720 11.250 ;
        RECT 39.670 6.900 40.300 11.250 ;
        RECT 41.260 6.900 41.890 11.250 ;
        RECT 42.830 6.900 43.460 11.250 ;
        RECT 43.790 8.050 44.480 10.470 ;
        RECT 44.740 6.890 45.370 11.240 ;
        RECT 46.330 6.890 46.960 11.240 ;
        RECT 47.900 6.900 48.530 11.250 ;
        RECT 49.480 6.900 50.110 11.250 ;
        RECT 51.070 6.900 51.700 11.250 ;
        RECT 52.640 6.900 53.270 11.250 ;
        RECT 54.550 6.920 55.180 11.270 ;
        RECT 56.140 6.920 56.770 11.270 ;
        RECT 57.710 6.930 58.340 11.280 ;
        RECT 59.290 6.930 59.920 11.280 ;
        RECT 60.880 6.930 61.510 11.280 ;
        RECT 62.450 6.930 63.080 11.280 ;
        RECT 63.350 8.010 64.040 10.430 ;
        RECT 64.340 6.920 64.970 11.270 ;
        RECT 65.930 6.920 66.560 11.270 ;
        RECT 67.500 6.930 68.130 11.280 ;
        RECT 69.080 6.930 69.710 11.280 ;
        RECT 70.670 6.930 71.300 11.280 ;
        RECT 72.240 6.930 72.870 11.280 ;
      LAYER met2 ;
        RECT 15.000 139.760 15.300 139.920 ;
        RECT 16.560 139.760 16.860 139.930 ;
        RECT 18.160 139.760 18.460 139.920 ;
        RECT 19.730 139.760 20.030 139.930 ;
        RECT 21.310 139.760 21.610 139.920 ;
        RECT 15.000 139.750 21.610 139.760 ;
        RECT 22.890 139.750 23.190 139.920 ;
        RECT 15.000 139.360 24.365 139.750 ;
        RECT 15.000 139.170 15.300 139.360 ;
        RECT 16.560 139.180 16.860 139.360 ;
        RECT 18.160 139.170 18.460 139.360 ;
        RECT 19.730 139.180 20.030 139.360 ;
        RECT 21.310 139.170 21.610 139.360 ;
        RECT 22.890 139.170 23.190 139.360 ;
        RECT 23.975 134.875 24.365 139.360 ;
        RECT 25.000 134.875 25.630 134.990 ;
        RECT 23.975 134.485 25.630 134.875 ;
        RECT 25.000 133.770 25.630 134.485 ;
        RECT 26.590 133.770 27.220 134.990 ;
        RECT 28.160 133.770 28.790 134.980 ;
        RECT 29.740 133.770 30.370 134.980 ;
        RECT 31.330 133.770 31.960 134.980 ;
        RECT 32.900 133.770 33.530 134.980 ;
        RECT 34.930 133.770 35.560 134.990 ;
        RECT 36.520 133.770 37.150 134.990 ;
        RECT 38.090 133.770 38.720 134.980 ;
        RECT 39.670 133.770 40.300 134.980 ;
        RECT 41.260 133.770 41.890 134.980 ;
        RECT 42.830 133.770 43.460 134.980 ;
        RECT 43.790 133.770 44.480 133.830 ;
        RECT 44.740 133.770 45.370 134.990 ;
        RECT 46.330 133.770 46.960 134.990 ;
        RECT 47.900 133.770 48.530 134.980 ;
        RECT 49.480 133.770 50.110 134.980 ;
        RECT 51.070 133.770 51.700 134.980 ;
        RECT 52.640 133.770 53.270 134.980 ;
        RECT 54.550 133.770 55.180 134.960 ;
        RECT 56.140 133.770 56.770 134.960 ;
        RECT 57.710 133.770 58.340 134.950 ;
        RECT 59.290 133.770 59.920 134.950 ;
        RECT 60.880 133.770 61.510 134.950 ;
        RECT 62.450 133.770 63.080 134.950 ;
        RECT 63.350 133.770 64.040 133.870 ;
        RECT 64.340 133.770 64.970 134.960 ;
        RECT 65.930 133.770 66.560 134.960 ;
        RECT 67.500 133.770 68.130 134.950 ;
        RECT 69.080 133.770 69.710 134.950 ;
        RECT 70.670 133.770 71.300 134.950 ;
        RECT 72.240 133.770 72.870 134.950 ;
        RECT 25.000 133.100 72.870 133.770 ;
        RECT 25.000 131.530 42.450 133.100 ;
        RECT 42.830 131.530 43.460 133.100 ;
        RECT 43.790 131.530 44.480 133.100 ;
        RECT 44.740 131.530 45.370 133.100 ;
        RECT 46.330 131.530 46.960 133.100 ;
        RECT 47.900 131.530 48.530 133.100 ;
        RECT 49.480 131.530 50.110 133.100 ;
        RECT 51.070 131.530 51.700 133.100 ;
        RECT 52.640 131.530 53.270 133.100 ;
        RECT 54.550 131.530 55.180 133.100 ;
        RECT 56.140 131.530 56.770 133.100 ;
        RECT 57.710 131.530 58.340 133.100 ;
        RECT 59.290 131.530 59.920 133.100 ;
        RECT 60.150 131.530 72.870 133.100 ;
        RECT 25.000 131.340 72.870 131.530 ;
        RECT 25.000 130.540 25.630 131.340 ;
        RECT 26.590 130.540 27.220 131.340 ;
        RECT 28.160 130.530 28.790 131.340 ;
        RECT 29.740 130.530 30.370 131.340 ;
        RECT 31.330 130.530 31.960 131.340 ;
        RECT 32.900 130.530 33.530 131.340 ;
        RECT 34.930 130.540 35.560 131.340 ;
        RECT 36.520 130.540 37.150 131.340 ;
        RECT 38.090 130.530 38.720 131.340 ;
        RECT 39.670 130.530 40.300 131.340 ;
        RECT 41.260 130.530 41.890 131.340 ;
        RECT 42.830 130.530 43.460 131.340 ;
        RECT 43.790 131.310 44.480 131.340 ;
        RECT 44.740 130.540 45.370 131.340 ;
        RECT 46.330 130.540 46.960 131.340 ;
        RECT 47.900 130.530 48.530 131.340 ;
        RECT 49.480 130.530 50.110 131.340 ;
        RECT 51.070 130.530 51.700 131.340 ;
        RECT 52.640 130.530 53.270 131.340 ;
        RECT 54.550 130.510 55.180 131.340 ;
        RECT 56.140 130.510 56.770 131.340 ;
        RECT 57.710 130.500 58.340 131.340 ;
        RECT 59.290 130.500 59.920 131.340 ;
        RECT 60.880 130.500 61.510 131.340 ;
        RECT 62.450 130.500 63.080 131.340 ;
        RECT 64.340 130.510 64.970 131.340 ;
        RECT 65.930 130.510 66.560 131.340 ;
        RECT 67.500 130.500 68.130 131.340 ;
        RECT 69.080 130.500 69.710 131.340 ;
        RECT 70.670 130.500 71.300 131.340 ;
        RECT 72.240 130.500 72.870 131.340 ;
        RECT 1.440 115.980 11.810 126.210 ;
        RECT 24.040 123.760 24.840 123.770 ;
        RECT 25.000 123.760 25.630 123.810 ;
        RECT 24.040 122.640 25.630 123.760 ;
        RECT 26.590 122.640 27.220 123.810 ;
        RECT 28.160 122.640 28.790 123.800 ;
        RECT 29.740 122.640 30.370 123.800 ;
        RECT 31.330 122.640 31.960 123.800 ;
        RECT 32.900 122.640 33.530 123.800 ;
        RECT 33.890 122.640 34.580 122.690 ;
        RECT 34.930 122.640 35.560 123.810 ;
        RECT 36.520 122.640 37.150 123.810 ;
        RECT 38.090 122.640 38.720 123.800 ;
        RECT 39.670 122.640 40.300 123.800 ;
        RECT 41.260 122.640 41.890 123.800 ;
        RECT 42.830 122.640 43.460 123.800 ;
        RECT 44.740 122.640 45.370 123.810 ;
        RECT 46.330 122.640 46.960 123.810 ;
        RECT 47.900 122.640 48.530 123.800 ;
        RECT 49.480 122.640 50.110 123.800 ;
        RECT 51.070 122.640 51.700 123.800 ;
        RECT 52.640 122.640 53.270 123.800 ;
        RECT 53.570 122.640 54.260 122.690 ;
        RECT 54.550 122.640 55.180 123.780 ;
        RECT 56.140 122.640 56.770 123.780 ;
        RECT 57.710 122.640 58.340 123.770 ;
        RECT 59.290 122.640 59.920 123.770 ;
        RECT 60.880 122.640 61.510 123.770 ;
        RECT 62.450 122.640 63.080 123.770 ;
        RECT 64.340 122.640 64.970 123.780 ;
        RECT 65.930 122.640 66.560 123.780 ;
        RECT 67.500 122.640 68.130 123.770 ;
        RECT 69.080 122.640 69.710 123.770 ;
        RECT 70.670 122.640 71.300 123.770 ;
        RECT 72.240 122.640 72.870 123.770 ;
        RECT 24.040 122.040 72.870 122.640 ;
        RECT 14.980 120.350 15.280 120.520 ;
        RECT 16.560 120.350 16.860 120.530 ;
        RECT 18.130 120.350 18.430 120.520 ;
        RECT 19.730 120.350 20.030 120.510 ;
        RECT 21.310 120.350 21.610 120.510 ;
        RECT 22.890 120.350 23.190 120.510 ;
        RECT 24.040 120.470 42.610 122.040 ;
        RECT 42.830 120.470 43.460 122.040 ;
        RECT 44.740 120.470 45.370 122.040 ;
        RECT 46.330 120.470 46.960 122.040 ;
        RECT 47.900 120.470 48.530 122.040 ;
        RECT 49.480 120.470 50.110 122.040 ;
        RECT 51.070 120.470 51.700 122.040 ;
        RECT 52.640 120.470 53.270 122.040 ;
        RECT 53.570 120.470 54.260 122.040 ;
        RECT 54.550 120.470 55.180 122.040 ;
        RECT 56.140 120.470 56.770 122.040 ;
        RECT 57.710 120.470 58.340 122.040 ;
        RECT 59.290 120.470 59.920 122.040 ;
        RECT 60.090 120.470 72.870 122.040 ;
        RECT 24.040 120.350 72.870 120.470 ;
        RECT 14.980 120.210 72.870 120.350 ;
        RECT 14.980 119.930 25.630 120.210 ;
        RECT 14.980 119.770 15.280 119.930 ;
        RECT 16.560 119.780 16.860 119.930 ;
        RECT 18.130 119.770 18.430 119.930 ;
        RECT 19.730 119.760 20.030 119.930 ;
        RECT 21.310 119.760 21.610 119.930 ;
        RECT 22.890 119.760 23.190 119.930 ;
        RECT 24.045 119.360 25.630 119.930 ;
        RECT 26.590 119.360 27.220 120.210 ;
        RECT 24.045 119.350 25.220 119.360 ;
        RECT 28.160 119.350 28.790 120.210 ;
        RECT 29.740 119.350 30.370 120.210 ;
        RECT 31.330 119.350 31.960 120.210 ;
        RECT 32.900 119.350 33.530 120.210 ;
        RECT 33.890 120.170 34.580 120.210 ;
        RECT 34.930 119.360 35.560 120.210 ;
        RECT 36.520 119.360 37.150 120.210 ;
        RECT 38.090 119.350 38.720 120.210 ;
        RECT 39.670 119.350 40.300 120.210 ;
        RECT 41.260 119.350 41.890 120.210 ;
        RECT 42.830 119.350 43.460 120.210 ;
        RECT 44.740 119.360 45.370 120.210 ;
        RECT 46.330 119.360 46.960 120.210 ;
        RECT 47.900 119.350 48.530 120.210 ;
        RECT 49.480 119.350 50.110 120.210 ;
        RECT 51.070 119.350 51.700 120.210 ;
        RECT 52.640 119.350 53.270 120.210 ;
        RECT 53.570 120.170 54.260 120.210 ;
        RECT 16.250 115.850 16.550 116.010 ;
        RECT 17.810 115.850 18.110 116.010 ;
        RECT 19.720 115.850 20.020 116.050 ;
        RECT 21.310 115.850 21.610 116.020 ;
        RECT 22.870 115.850 23.170 116.020 ;
        RECT 24.045 115.850 24.435 119.350 ;
        RECT 54.550 119.330 55.180 120.210 ;
        RECT 56.140 119.330 56.770 120.210 ;
        RECT 57.710 119.320 58.340 120.210 ;
        RECT 59.290 119.320 59.920 120.210 ;
        RECT 60.880 119.320 61.510 120.210 ;
        RECT 62.450 119.320 63.080 120.210 ;
        RECT 64.340 119.330 64.970 120.210 ;
        RECT 65.930 119.330 66.560 120.210 ;
        RECT 67.500 119.320 68.130 120.210 ;
        RECT 69.080 119.320 69.710 120.210 ;
        RECT 70.670 119.320 71.300 120.210 ;
        RECT 72.240 119.320 72.870 120.210 ;
        RECT 16.250 115.460 24.435 115.850 ;
        RECT 16.250 115.260 16.550 115.460 ;
        RECT 17.810 115.260 18.110 115.460 ;
        RECT 18.605 111.195 18.995 115.460 ;
        RECT 19.720 115.300 20.020 115.460 ;
        RECT 21.310 115.270 21.610 115.460 ;
        RECT 22.870 115.270 23.170 115.460 ;
        RECT 16.975 110.805 18.995 111.195 ;
        RECT 25.000 111.380 25.630 112.630 ;
        RECT 26.590 111.380 27.220 112.630 ;
        RECT 28.160 111.380 28.790 112.620 ;
        RECT 29.740 111.380 30.370 112.620 ;
        RECT 31.330 111.380 31.960 112.620 ;
        RECT 32.900 111.380 33.530 112.620 ;
        RECT 34.930 111.380 35.560 112.630 ;
        RECT 36.520 111.380 37.150 112.630 ;
        RECT 38.090 111.380 38.720 112.620 ;
        RECT 39.670 111.380 40.300 112.620 ;
        RECT 41.260 111.380 41.890 112.620 ;
        RECT 42.830 111.380 43.460 112.620 ;
        RECT 43.780 111.380 44.470 111.440 ;
        RECT 44.740 111.380 45.370 112.630 ;
        RECT 46.330 111.380 46.960 112.630 ;
        RECT 47.900 111.380 48.530 112.620 ;
        RECT 49.480 111.380 50.110 112.620 ;
        RECT 51.070 111.380 51.700 112.620 ;
        RECT 52.640 111.380 53.270 112.620 ;
        RECT 54.550 111.380 55.180 112.600 ;
        RECT 56.140 111.380 56.770 112.600 ;
        RECT 57.710 111.380 58.340 112.590 ;
        RECT 59.290 111.380 59.920 112.590 ;
        RECT 60.880 111.380 61.510 112.590 ;
        RECT 62.450 111.380 63.080 112.590 ;
        RECT 63.360 111.380 64.050 111.420 ;
        RECT 64.340 111.380 64.970 112.600 ;
        RECT 65.930 111.380 66.560 112.600 ;
        RECT 67.500 111.380 68.130 112.590 ;
        RECT 69.080 111.380 69.710 112.590 ;
        RECT 70.670 111.380 71.300 112.590 ;
        RECT 72.240 111.380 72.870 112.590 ;
        RECT 16.975 109.135 17.365 110.805 ;
        RECT 25.000 110.770 72.870 111.380 ;
        RECT 25.000 109.200 42.520 110.770 ;
        RECT 42.830 109.200 43.460 110.770 ;
        RECT 43.780 109.200 44.470 110.770 ;
        RECT 44.740 109.200 45.370 110.770 ;
        RECT 46.330 109.200 46.960 110.770 ;
        RECT 47.900 109.200 48.530 110.770 ;
        RECT 49.480 109.200 50.110 110.770 ;
        RECT 51.070 109.200 51.700 110.770 ;
        RECT 52.640 109.200 53.270 110.770 ;
        RECT 54.550 109.200 55.180 110.770 ;
        RECT 56.140 109.200 56.770 110.770 ;
        RECT 57.710 109.200 58.340 110.770 ;
        RECT 59.290 109.200 59.920 110.770 ;
        RECT 60.120 109.200 72.870 110.770 ;
        RECT 25.000 108.950 72.870 109.200 ;
        RECT 25.000 108.180 25.630 108.950 ;
        RECT 26.590 108.180 27.220 108.950 ;
        RECT 28.160 108.170 28.790 108.950 ;
        RECT 29.740 108.170 30.370 108.950 ;
        RECT 31.330 108.170 31.960 108.950 ;
        RECT 32.900 108.170 33.530 108.950 ;
        RECT 34.930 108.180 35.560 108.950 ;
        RECT 36.520 108.180 37.150 108.950 ;
        RECT 38.090 108.170 38.720 108.950 ;
        RECT 39.670 108.170 40.300 108.950 ;
        RECT 41.260 108.170 41.890 108.950 ;
        RECT 42.830 108.170 43.460 108.950 ;
        RECT 43.780 108.920 44.470 108.950 ;
        RECT 44.740 108.180 45.370 108.950 ;
        RECT 46.330 108.180 46.960 108.950 ;
        RECT 47.900 108.170 48.530 108.950 ;
        RECT 49.480 108.170 50.110 108.950 ;
        RECT 51.070 108.170 51.700 108.950 ;
        RECT 52.640 108.170 53.270 108.950 ;
        RECT 54.550 108.150 55.180 108.950 ;
        RECT 56.140 108.150 56.770 108.950 ;
        RECT 57.710 108.140 58.340 108.950 ;
        RECT 59.290 108.140 59.920 108.950 ;
        RECT 60.880 108.140 61.510 108.950 ;
        RECT 62.450 108.140 63.080 108.950 ;
        RECT 63.360 108.900 64.050 108.950 ;
        RECT 64.340 108.150 64.970 108.950 ;
        RECT 65.930 108.150 66.560 108.950 ;
        RECT 67.500 108.140 68.130 108.950 ;
        RECT 69.080 108.140 69.710 108.950 ;
        RECT 70.670 108.140 71.300 108.950 ;
        RECT 72.240 108.140 72.870 108.950 ;
        RECT 25.000 100.430 25.630 101.450 ;
        RECT 26.590 100.430 27.220 101.450 ;
        RECT 28.160 100.430 28.790 101.440 ;
        RECT 29.740 100.430 30.370 101.440 ;
        RECT 31.330 100.430 31.960 101.440 ;
        RECT 32.900 100.430 33.530 101.440 ;
        RECT 33.870 100.430 34.560 100.500 ;
        RECT 34.930 100.430 35.560 101.450 ;
        RECT 36.520 100.430 37.150 101.450 ;
        RECT 38.090 100.430 38.720 101.440 ;
        RECT 39.670 100.430 40.300 101.440 ;
        RECT 41.260 100.430 41.890 101.440 ;
        RECT 42.830 100.430 43.460 101.440 ;
        RECT 44.740 100.430 45.370 101.450 ;
        RECT 46.330 100.430 46.960 101.450 ;
        RECT 47.900 100.430 48.530 101.440 ;
        RECT 49.480 100.430 50.110 101.440 ;
        RECT 51.070 100.430 51.700 101.440 ;
        RECT 52.640 100.430 53.270 101.440 ;
        RECT 53.600 100.430 54.290 100.460 ;
        RECT 54.550 100.430 55.180 101.420 ;
        RECT 56.140 100.430 56.770 101.420 ;
        RECT 57.710 100.430 58.340 101.410 ;
        RECT 59.290 100.430 59.920 101.410 ;
        RECT 60.880 100.430 61.510 101.410 ;
        RECT 62.450 100.430 63.080 101.410 ;
        RECT 64.340 100.430 64.970 101.420 ;
        RECT 65.930 100.430 66.560 101.420 ;
        RECT 67.500 100.430 68.130 101.410 ;
        RECT 69.080 100.430 69.710 101.410 ;
        RECT 70.670 100.430 71.300 101.410 ;
        RECT 72.240 100.430 72.870 101.410 ;
        RECT 25.000 100.160 72.870 100.430 ;
        RECT 25.000 98.590 42.665 100.160 ;
        RECT 42.830 98.590 43.460 100.160 ;
        RECT 44.740 98.590 45.370 100.160 ;
        RECT 46.330 98.590 46.960 100.160 ;
        RECT 47.900 98.590 48.530 100.160 ;
        RECT 49.480 98.590 50.110 100.160 ;
        RECT 51.070 98.590 51.700 100.160 ;
        RECT 52.640 98.590 53.270 100.160 ;
        RECT 53.600 98.590 54.290 100.160 ;
        RECT 54.550 98.590 55.180 100.160 ;
        RECT 56.140 98.590 56.770 100.160 ;
        RECT 57.710 98.590 58.340 100.160 ;
        RECT 59.290 98.590 59.920 100.160 ;
        RECT 60.150 98.590 72.870 100.160 ;
        RECT 25.000 98.000 72.870 98.590 ;
        RECT 25.000 97.000 25.630 98.000 ;
        RECT 26.590 97.000 27.220 98.000 ;
        RECT 28.160 96.990 28.790 98.000 ;
        RECT 29.740 96.990 30.370 98.000 ;
        RECT 31.330 96.990 31.960 98.000 ;
        RECT 32.900 96.990 33.530 98.000 ;
        RECT 33.870 97.980 34.560 98.000 ;
        RECT 34.930 97.000 35.560 98.000 ;
        RECT 36.520 97.000 37.150 98.000 ;
        RECT 38.090 96.990 38.720 98.000 ;
        RECT 39.670 96.990 40.300 98.000 ;
        RECT 41.260 96.990 41.890 98.000 ;
        RECT 42.830 96.990 43.460 98.000 ;
        RECT 44.740 97.000 45.370 98.000 ;
        RECT 46.330 97.000 46.960 98.000 ;
        RECT 47.900 96.990 48.530 98.000 ;
        RECT 49.480 96.990 50.110 98.000 ;
        RECT 51.070 96.990 51.700 98.000 ;
        RECT 52.640 96.990 53.270 98.000 ;
        RECT 53.600 97.940 54.290 98.000 ;
        RECT 54.550 96.970 55.180 98.000 ;
        RECT 56.140 96.970 56.770 98.000 ;
        RECT 57.710 96.960 58.340 98.000 ;
        RECT 59.290 96.960 59.920 98.000 ;
        RECT 60.880 96.960 61.510 98.000 ;
        RECT 62.450 96.960 63.080 98.000 ;
        RECT 64.340 96.970 64.970 98.000 ;
        RECT 65.930 96.970 66.560 98.000 ;
        RECT 67.500 96.960 68.130 98.000 ;
        RECT 69.080 96.960 69.710 98.000 ;
        RECT 70.670 96.960 71.300 98.000 ;
        RECT 72.240 96.960 72.870 98.000 ;
        RECT 3.305 80.455 3.595 80.505 ;
        RECT 4.885 80.455 5.175 80.505 ;
        RECT 6.465 80.455 6.755 80.505 ;
        RECT 7.935 80.455 8.205 80.505 ;
        RECT 9.385 80.455 9.675 80.505 ;
        RECT 10.965 80.455 11.255 80.505 ;
        RECT 12.545 80.455 12.835 80.505 ;
        RECT 3.305 80.285 13.155 80.455 ;
        RECT 3.305 80.280 13.710 80.285 ;
        RECT 3.305 79.875 14.260 80.280 ;
        RECT 3.305 79.855 13.155 79.875 ;
        RECT 3.305 79.805 3.595 79.855 ;
        RECT 4.885 79.805 5.175 79.855 ;
        RECT 6.465 79.805 6.755 79.855 ;
        RECT 7.935 79.805 8.205 79.855 ;
        RECT 9.385 79.805 9.675 79.855 ;
        RECT 10.965 79.805 11.255 79.855 ;
        RECT 12.545 79.805 12.835 79.855 ;
        RECT 13.710 79.585 14.260 79.875 ;
        RECT 17.695 79.800 17.955 79.850 ;
        RECT 19.275 79.800 19.535 79.850 ;
        RECT 19.945 79.800 20.365 79.850 ;
        RECT 20.775 79.800 21.035 79.850 ;
        RECT 22.355 79.800 22.615 79.850 ;
        RECT 22.975 79.800 23.825 79.845 ;
        RECT 17.695 79.585 23.825 79.800 ;
        RECT 13.710 79.180 23.825 79.585 ;
        RECT 14.260 79.175 23.825 79.180 ;
        RECT 17.695 78.950 23.825 79.175 ;
        RECT 17.695 78.900 17.955 78.950 ;
        RECT 19.275 78.900 19.535 78.950 ;
        RECT 19.945 78.900 20.365 78.950 ;
        RECT 20.775 78.900 21.035 78.950 ;
        RECT 22.355 78.900 22.615 78.950 ;
        RECT 22.975 78.905 23.825 78.950 ;
        RECT 25.000 43.830 25.630 44.830 ;
        RECT 26.590 43.830 27.220 44.830 ;
        RECT 28.160 43.830 28.790 44.840 ;
        RECT 29.740 43.830 30.370 44.840 ;
        RECT 31.330 43.830 31.960 44.840 ;
        RECT 32.900 43.830 33.530 44.840 ;
        RECT 33.870 43.830 34.560 43.850 ;
        RECT 34.930 43.830 35.560 44.830 ;
        RECT 36.520 43.830 37.150 44.830 ;
        RECT 38.090 43.830 38.720 44.840 ;
        RECT 39.670 43.830 40.300 44.840 ;
        RECT 41.260 43.830 41.890 44.840 ;
        RECT 42.830 43.830 43.460 44.840 ;
        RECT 44.740 43.830 45.370 44.830 ;
        RECT 46.330 43.830 46.960 44.830 ;
        RECT 47.900 43.830 48.530 44.840 ;
        RECT 49.480 43.830 50.110 44.840 ;
        RECT 51.070 43.830 51.700 44.840 ;
        RECT 52.640 43.830 53.270 44.840 ;
        RECT 53.600 43.830 54.290 43.890 ;
        RECT 54.550 43.830 55.180 44.860 ;
        RECT 56.140 43.830 56.770 44.860 ;
        RECT 57.710 43.830 58.340 44.870 ;
        RECT 59.290 43.830 59.920 44.870 ;
        RECT 60.880 43.830 61.510 44.870 ;
        RECT 62.450 43.830 63.080 44.870 ;
        RECT 64.340 43.830 64.970 44.860 ;
        RECT 65.930 43.830 66.560 44.860 ;
        RECT 67.500 43.830 68.130 44.870 ;
        RECT 69.080 43.830 69.710 44.870 ;
        RECT 70.670 43.830 71.300 44.870 ;
        RECT 72.240 43.830 72.870 44.870 ;
        RECT 25.000 43.240 72.870 43.830 ;
        RECT 25.000 41.670 42.665 43.240 ;
        RECT 42.830 41.670 43.460 43.240 ;
        RECT 44.740 41.670 45.370 43.240 ;
        RECT 46.330 41.670 46.960 43.240 ;
        RECT 47.900 41.670 48.530 43.240 ;
        RECT 49.480 41.670 50.110 43.240 ;
        RECT 51.070 41.670 51.700 43.240 ;
        RECT 52.640 41.670 53.270 43.240 ;
        RECT 53.600 41.670 54.290 43.240 ;
        RECT 54.550 41.670 55.180 43.240 ;
        RECT 56.140 41.670 56.770 43.240 ;
        RECT 57.710 41.670 58.340 43.240 ;
        RECT 59.290 41.670 59.920 43.240 ;
        RECT 60.150 41.670 72.870 43.240 ;
        RECT 25.000 41.400 72.870 41.670 ;
        RECT 25.000 40.380 25.630 41.400 ;
        RECT 26.590 40.380 27.220 41.400 ;
        RECT 28.160 40.390 28.790 41.400 ;
        RECT 29.740 40.390 30.370 41.400 ;
        RECT 31.330 40.390 31.960 41.400 ;
        RECT 32.900 40.390 33.530 41.400 ;
        RECT 33.870 41.330 34.560 41.400 ;
        RECT 34.930 40.380 35.560 41.400 ;
        RECT 36.520 40.380 37.150 41.400 ;
        RECT 38.090 40.390 38.720 41.400 ;
        RECT 39.670 40.390 40.300 41.400 ;
        RECT 41.260 40.390 41.890 41.400 ;
        RECT 42.830 40.390 43.460 41.400 ;
        RECT 44.740 40.380 45.370 41.400 ;
        RECT 46.330 40.380 46.960 41.400 ;
        RECT 47.900 40.390 48.530 41.400 ;
        RECT 49.480 40.390 50.110 41.400 ;
        RECT 51.070 40.390 51.700 41.400 ;
        RECT 52.640 40.390 53.270 41.400 ;
        RECT 53.600 41.370 54.290 41.400 ;
        RECT 54.550 40.410 55.180 41.400 ;
        RECT 56.140 40.410 56.770 41.400 ;
        RECT 57.710 40.420 58.340 41.400 ;
        RECT 59.290 40.420 59.920 41.400 ;
        RECT 60.880 40.420 61.510 41.400 ;
        RECT 62.450 40.420 63.080 41.400 ;
        RECT 64.340 40.410 64.970 41.400 ;
        RECT 65.930 40.410 66.560 41.400 ;
        RECT 67.500 40.420 68.130 41.400 ;
        RECT 69.080 40.420 69.710 41.400 ;
        RECT 70.670 40.420 71.300 41.400 ;
        RECT 72.240 40.420 72.870 41.400 ;
        RECT 25.000 32.880 25.630 33.650 ;
        RECT 26.590 32.880 27.220 33.650 ;
        RECT 28.160 32.880 28.790 33.660 ;
        RECT 29.740 32.880 30.370 33.660 ;
        RECT 31.330 32.880 31.960 33.660 ;
        RECT 32.900 32.880 33.530 33.660 ;
        RECT 34.930 32.880 35.560 33.650 ;
        RECT 36.520 32.880 37.150 33.650 ;
        RECT 38.090 32.880 38.720 33.660 ;
        RECT 39.670 32.880 40.300 33.660 ;
        RECT 41.260 32.880 41.890 33.660 ;
        RECT 42.830 32.880 43.460 33.660 ;
        RECT 43.780 32.880 44.470 32.910 ;
        RECT 44.740 32.880 45.370 33.650 ;
        RECT 46.330 32.880 46.960 33.650 ;
        RECT 47.900 32.880 48.530 33.660 ;
        RECT 49.480 32.880 50.110 33.660 ;
        RECT 51.070 32.880 51.700 33.660 ;
        RECT 52.640 32.880 53.270 33.660 ;
        RECT 54.550 32.880 55.180 33.680 ;
        RECT 56.140 32.880 56.770 33.680 ;
        RECT 57.710 32.880 58.340 33.690 ;
        RECT 59.290 32.880 59.920 33.690 ;
        RECT 60.880 32.880 61.510 33.690 ;
        RECT 62.450 32.880 63.080 33.690 ;
        RECT 63.360 32.880 64.050 32.930 ;
        RECT 64.340 32.880 64.970 33.680 ;
        RECT 65.930 32.880 66.560 33.680 ;
        RECT 67.500 32.880 68.130 33.690 ;
        RECT 69.080 32.880 69.710 33.690 ;
        RECT 70.670 32.880 71.300 33.690 ;
        RECT 72.240 32.880 72.870 33.690 ;
        RECT 16.975 31.025 17.365 32.695 ;
        RECT 25.000 32.630 72.870 32.880 ;
        RECT 25.000 31.060 42.520 32.630 ;
        RECT 42.830 31.060 43.460 32.630 ;
        RECT 43.780 31.060 44.470 32.630 ;
        RECT 44.740 31.060 45.370 32.630 ;
        RECT 46.330 31.060 46.960 32.630 ;
        RECT 47.900 31.060 48.530 32.630 ;
        RECT 49.480 31.060 50.110 32.630 ;
        RECT 51.070 31.060 51.700 32.630 ;
        RECT 52.640 31.060 53.270 32.630 ;
        RECT 54.550 31.060 55.180 32.630 ;
        RECT 56.140 31.060 56.770 32.630 ;
        RECT 57.710 31.060 58.340 32.630 ;
        RECT 59.290 31.060 59.920 32.630 ;
        RECT 60.120 31.060 72.870 32.630 ;
        RECT 16.975 30.635 18.995 31.025 ;
        RECT 1.300 18.350 11.780 28.310 ;
        RECT 16.250 26.370 16.550 26.570 ;
        RECT 17.810 26.370 18.110 26.570 ;
        RECT 18.605 26.370 18.995 30.635 ;
        RECT 25.000 30.450 72.870 31.060 ;
        RECT 25.000 29.200 25.630 30.450 ;
        RECT 26.590 29.200 27.220 30.450 ;
        RECT 28.160 29.210 28.790 30.450 ;
        RECT 29.740 29.210 30.370 30.450 ;
        RECT 31.330 29.210 31.960 30.450 ;
        RECT 32.900 29.210 33.530 30.450 ;
        RECT 34.930 29.200 35.560 30.450 ;
        RECT 36.520 29.200 37.150 30.450 ;
        RECT 38.090 29.210 38.720 30.450 ;
        RECT 39.670 29.210 40.300 30.450 ;
        RECT 41.260 29.210 41.890 30.450 ;
        RECT 42.830 29.210 43.460 30.450 ;
        RECT 43.780 30.390 44.470 30.450 ;
        RECT 44.740 29.200 45.370 30.450 ;
        RECT 46.330 29.200 46.960 30.450 ;
        RECT 47.900 29.210 48.530 30.450 ;
        RECT 49.480 29.210 50.110 30.450 ;
        RECT 51.070 29.210 51.700 30.450 ;
        RECT 52.640 29.210 53.270 30.450 ;
        RECT 54.550 29.230 55.180 30.450 ;
        RECT 56.140 29.230 56.770 30.450 ;
        RECT 57.710 29.240 58.340 30.450 ;
        RECT 59.290 29.240 59.920 30.450 ;
        RECT 60.880 29.240 61.510 30.450 ;
        RECT 62.450 29.240 63.080 30.450 ;
        RECT 63.360 30.410 64.050 30.450 ;
        RECT 64.340 29.230 64.970 30.450 ;
        RECT 65.930 29.230 66.560 30.450 ;
        RECT 67.500 29.240 68.130 30.450 ;
        RECT 69.080 29.240 69.710 30.450 ;
        RECT 70.670 29.240 71.300 30.450 ;
        RECT 72.240 29.240 72.870 30.450 ;
        RECT 19.720 26.370 20.020 26.530 ;
        RECT 21.310 26.370 21.610 26.560 ;
        RECT 22.870 26.370 23.170 26.560 ;
        RECT 16.250 25.980 24.435 26.370 ;
        RECT 16.250 25.820 16.550 25.980 ;
        RECT 17.810 25.820 18.110 25.980 ;
        RECT 19.720 25.780 20.020 25.980 ;
        RECT 21.310 25.810 21.610 25.980 ;
        RECT 22.870 25.810 23.170 25.980 ;
        RECT 24.045 22.480 24.435 25.980 ;
        RECT 24.045 22.470 25.220 22.480 ;
        RECT 14.980 21.900 15.280 22.060 ;
        RECT 16.560 21.900 16.860 22.050 ;
        RECT 18.130 21.900 18.430 22.060 ;
        RECT 19.730 21.900 20.030 22.070 ;
        RECT 21.310 21.900 21.610 22.070 ;
        RECT 22.890 21.900 23.190 22.070 ;
        RECT 24.045 21.900 25.630 22.470 ;
        RECT 14.980 21.620 25.630 21.900 ;
        RECT 26.590 21.620 27.220 22.470 ;
        RECT 28.160 21.620 28.790 22.480 ;
        RECT 29.740 21.620 30.370 22.480 ;
        RECT 31.330 21.620 31.960 22.480 ;
        RECT 32.900 21.620 33.530 22.480 ;
        RECT 33.890 21.620 34.580 21.660 ;
        RECT 34.930 21.620 35.560 22.470 ;
        RECT 36.520 21.620 37.150 22.470 ;
        RECT 38.090 21.620 38.720 22.480 ;
        RECT 39.670 21.620 40.300 22.480 ;
        RECT 41.260 21.620 41.890 22.480 ;
        RECT 42.830 21.620 43.460 22.480 ;
        RECT 44.740 21.620 45.370 22.470 ;
        RECT 46.330 21.620 46.960 22.470 ;
        RECT 47.900 21.620 48.530 22.480 ;
        RECT 49.480 21.620 50.110 22.480 ;
        RECT 51.070 21.620 51.700 22.480 ;
        RECT 52.640 21.620 53.270 22.480 ;
        RECT 53.570 21.620 54.260 21.660 ;
        RECT 54.550 21.620 55.180 22.500 ;
        RECT 56.140 21.620 56.770 22.500 ;
        RECT 57.710 21.620 58.340 22.510 ;
        RECT 59.290 21.620 59.920 22.510 ;
        RECT 60.880 21.620 61.510 22.510 ;
        RECT 62.450 21.620 63.080 22.510 ;
        RECT 64.340 21.620 64.970 22.500 ;
        RECT 65.930 21.620 66.560 22.500 ;
        RECT 67.500 21.620 68.130 22.510 ;
        RECT 69.080 21.620 69.710 22.510 ;
        RECT 70.670 21.620 71.300 22.510 ;
        RECT 72.240 21.620 72.870 22.510 ;
        RECT 14.980 21.480 72.870 21.620 ;
        RECT 14.980 21.310 15.280 21.480 ;
        RECT 16.560 21.300 16.860 21.480 ;
        RECT 18.130 21.310 18.430 21.480 ;
        RECT 19.730 21.320 20.030 21.480 ;
        RECT 21.310 21.320 21.610 21.480 ;
        RECT 22.890 21.320 23.190 21.480 ;
        RECT 24.040 21.360 72.870 21.480 ;
        RECT 24.040 19.790 42.610 21.360 ;
        RECT 42.830 19.790 43.460 21.360 ;
        RECT 44.740 19.790 45.370 21.360 ;
        RECT 46.330 19.790 46.960 21.360 ;
        RECT 47.900 19.790 48.530 21.360 ;
        RECT 49.480 19.790 50.110 21.360 ;
        RECT 51.070 19.790 51.700 21.360 ;
        RECT 52.640 19.790 53.270 21.360 ;
        RECT 53.570 19.790 54.260 21.360 ;
        RECT 54.550 19.790 55.180 21.360 ;
        RECT 56.140 19.790 56.770 21.360 ;
        RECT 57.710 19.790 58.340 21.360 ;
        RECT 59.290 19.790 59.920 21.360 ;
        RECT 60.090 19.790 72.870 21.360 ;
        RECT 24.040 19.190 72.870 19.790 ;
        RECT 24.040 18.070 25.630 19.190 ;
        RECT 24.040 18.060 24.840 18.070 ;
        RECT 25.000 18.020 25.630 18.070 ;
        RECT 26.590 18.020 27.220 19.190 ;
        RECT 28.160 18.030 28.790 19.190 ;
        RECT 29.740 18.030 30.370 19.190 ;
        RECT 31.330 18.030 31.960 19.190 ;
        RECT 32.900 18.030 33.530 19.190 ;
        RECT 33.890 19.140 34.580 19.190 ;
        RECT 34.930 18.020 35.560 19.190 ;
        RECT 36.520 18.020 37.150 19.190 ;
        RECT 38.090 18.030 38.720 19.190 ;
        RECT 39.670 18.030 40.300 19.190 ;
        RECT 41.260 18.030 41.890 19.190 ;
        RECT 42.830 18.030 43.460 19.190 ;
        RECT 44.740 18.020 45.370 19.190 ;
        RECT 46.330 18.020 46.960 19.190 ;
        RECT 47.900 18.030 48.530 19.190 ;
        RECT 49.480 18.030 50.110 19.190 ;
        RECT 51.070 18.030 51.700 19.190 ;
        RECT 52.640 18.030 53.270 19.190 ;
        RECT 53.570 19.140 54.260 19.190 ;
        RECT 54.550 18.050 55.180 19.190 ;
        RECT 56.140 18.050 56.770 19.190 ;
        RECT 57.710 18.060 58.340 19.190 ;
        RECT 59.290 18.060 59.920 19.190 ;
        RECT 60.880 18.060 61.510 19.190 ;
        RECT 62.450 18.060 63.080 19.190 ;
        RECT 64.340 18.050 64.970 19.190 ;
        RECT 65.930 18.050 66.560 19.190 ;
        RECT 67.500 18.060 68.130 19.190 ;
        RECT 69.080 18.060 69.710 19.190 ;
        RECT 70.670 18.060 71.300 19.190 ;
        RECT 72.240 18.060 72.870 19.190 ;
        RECT 25.000 10.490 25.630 11.290 ;
        RECT 26.590 10.490 27.220 11.290 ;
        RECT 28.160 10.490 28.790 11.300 ;
        RECT 29.740 10.490 30.370 11.300 ;
        RECT 31.330 10.490 31.960 11.300 ;
        RECT 32.900 10.490 33.530 11.300 ;
        RECT 34.930 10.490 35.560 11.290 ;
        RECT 36.520 10.490 37.150 11.290 ;
        RECT 38.090 10.490 38.720 11.300 ;
        RECT 39.670 10.490 40.300 11.300 ;
        RECT 41.260 10.490 41.890 11.300 ;
        RECT 42.830 10.490 43.460 11.300 ;
        RECT 43.790 10.490 44.480 10.520 ;
        RECT 44.740 10.490 45.370 11.290 ;
        RECT 46.330 10.490 46.960 11.290 ;
        RECT 47.900 10.490 48.530 11.300 ;
        RECT 49.480 10.490 50.110 11.300 ;
        RECT 51.070 10.490 51.700 11.300 ;
        RECT 52.640 10.490 53.270 11.300 ;
        RECT 54.550 10.490 55.180 11.320 ;
        RECT 56.140 10.490 56.770 11.320 ;
        RECT 57.710 10.490 58.340 11.330 ;
        RECT 59.290 10.490 59.920 11.330 ;
        RECT 60.880 10.490 61.510 11.330 ;
        RECT 62.450 10.490 63.080 11.330 ;
        RECT 64.340 10.490 64.970 11.320 ;
        RECT 65.930 10.490 66.560 11.320 ;
        RECT 67.500 10.490 68.130 11.330 ;
        RECT 69.080 10.490 69.710 11.330 ;
        RECT 70.670 10.490 71.300 11.330 ;
        RECT 72.240 10.490 72.870 11.330 ;
        RECT 25.000 10.300 72.870 10.490 ;
        RECT 25.000 8.730 42.450 10.300 ;
        RECT 42.830 8.730 43.460 10.300 ;
        RECT 43.790 8.730 44.480 10.300 ;
        RECT 44.740 8.730 45.370 10.300 ;
        RECT 46.330 8.730 46.960 10.300 ;
        RECT 47.900 8.730 48.530 10.300 ;
        RECT 49.480 8.730 50.110 10.300 ;
        RECT 51.070 8.730 51.700 10.300 ;
        RECT 52.640 8.730 53.270 10.300 ;
        RECT 54.550 8.730 55.180 10.300 ;
        RECT 56.140 8.730 56.770 10.300 ;
        RECT 57.710 8.730 58.340 10.300 ;
        RECT 59.290 8.730 59.920 10.300 ;
        RECT 60.150 8.730 72.870 10.300 ;
        RECT 25.000 8.060 72.870 8.730 ;
        RECT 25.000 7.345 25.630 8.060 ;
        RECT 23.975 6.955 25.630 7.345 ;
        RECT 15.000 2.470 15.300 2.660 ;
        RECT 16.560 2.470 16.860 2.650 ;
        RECT 18.160 2.470 18.460 2.660 ;
        RECT 19.730 2.470 20.030 2.650 ;
        RECT 21.310 2.470 21.610 2.660 ;
        RECT 22.890 2.470 23.190 2.660 ;
        RECT 23.975 2.470 24.365 6.955 ;
        RECT 25.000 6.840 25.630 6.955 ;
        RECT 26.590 6.840 27.220 8.060 ;
        RECT 28.160 6.850 28.790 8.060 ;
        RECT 29.740 6.850 30.370 8.060 ;
        RECT 31.330 6.850 31.960 8.060 ;
        RECT 32.900 6.850 33.530 8.060 ;
        RECT 34.930 6.840 35.560 8.060 ;
        RECT 36.520 6.840 37.150 8.060 ;
        RECT 38.090 6.850 38.720 8.060 ;
        RECT 39.670 6.850 40.300 8.060 ;
        RECT 41.260 6.850 41.890 8.060 ;
        RECT 42.830 6.850 43.460 8.060 ;
        RECT 43.790 8.000 44.480 8.060 ;
        RECT 44.740 6.840 45.370 8.060 ;
        RECT 46.330 6.840 46.960 8.060 ;
        RECT 47.900 6.850 48.530 8.060 ;
        RECT 49.480 6.850 50.110 8.060 ;
        RECT 51.070 6.850 51.700 8.060 ;
        RECT 52.640 6.850 53.270 8.060 ;
        RECT 54.550 6.870 55.180 8.060 ;
        RECT 56.140 6.870 56.770 8.060 ;
        RECT 57.710 6.880 58.340 8.060 ;
        RECT 59.290 6.880 59.920 8.060 ;
        RECT 60.880 6.880 61.510 8.060 ;
        RECT 62.450 6.880 63.080 8.060 ;
        RECT 63.350 7.960 64.040 8.060 ;
        RECT 64.340 6.870 64.970 8.060 ;
        RECT 65.930 6.870 66.560 8.060 ;
        RECT 67.500 6.880 68.130 8.060 ;
        RECT 69.080 6.880 69.710 8.060 ;
        RECT 70.670 6.880 71.300 8.060 ;
        RECT 72.240 6.880 72.870 8.060 ;
        RECT 15.000 2.080 24.365 2.470 ;
        RECT 15.000 2.070 21.610 2.080 ;
        RECT 15.000 1.910 15.300 2.070 ;
        RECT 16.560 1.900 16.860 2.070 ;
        RECT 18.160 1.910 18.460 2.070 ;
        RECT 19.730 1.900 20.030 2.070 ;
        RECT 21.310 1.910 21.610 2.070 ;
        RECT 22.890 1.910 23.190 2.080 ;
      LAYER via2 ;
        RECT 27.480 131.530 42.450 133.100 ;
        RECT 1.440 116.030 11.810 126.160 ;
        RECT 27.420 120.470 42.610 122.040 ;
        RECT 27.450 109.200 42.520 110.770 ;
        RECT 27.480 98.590 42.665 100.160 ;
        RECT 22.975 78.950 23.825 79.800 ;
        RECT 27.480 41.670 42.665 43.240 ;
        RECT 27.450 31.060 42.520 32.630 ;
        RECT 1.300 18.400 11.780 28.260 ;
        RECT 27.420 19.790 42.610 21.360 ;
        RECT 27.480 8.730 42.450 10.300 ;
      LAYER met3 ;
        RECT 27.270 126.300 42.690 133.380 ;
        RECT 1.440 126.185 42.690 126.300 ;
        RECT 1.390 116.030 42.690 126.185 ;
        RECT 1.390 116.005 11.860 116.030 ;
        RECT 27.270 79.830 42.690 116.030 ;
        RECT 22.920 78.900 42.690 79.830 ;
        RECT 27.270 28.310 42.690 78.900 ;
        RECT 1.250 18.380 42.690 28.310 ;
        RECT 1.250 18.375 11.830 18.380 ;
        RECT 27.270 8.450 42.690 18.380 ;
      LAYER via3 ;
        RECT 27.490 75.500 42.300 98.250 ;
      LAYER met4 ;
        RECT 0.460 134.660 72.360 141.240 ;
        RECT 0.350 129.230 73.700 134.660 ;
        RECT 0.460 75.220 72.360 129.230 ;
      LAYER met5 ;
        RECT 0.230 129.110 73.820 134.780 ;
    END
  END vdd
  PIN in_hi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 90.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.245 75.505 2.145 75.675 ;
        RECT 2.435 75.505 3.335 75.675 ;
        RECT 3.625 75.505 4.525 75.675 ;
        RECT 4.815 75.505 5.715 75.675 ;
        RECT 6.005 75.505 6.905 75.675 ;
        RECT 9.095 75.505 9.995 75.675 ;
        RECT 10.285 75.505 11.185 75.675 ;
        RECT 11.475 75.505 12.375 75.675 ;
        RECT 12.665 75.505 13.565 75.675 ;
        RECT 13.855 75.505 14.755 75.675 ;
        RECT 1.245 64.955 2.145 65.125 ;
        RECT 2.435 64.955 3.335 65.125 ;
        RECT 3.625 64.955 4.525 65.125 ;
        RECT 4.815 64.955 5.715 65.125 ;
        RECT 6.005 64.955 6.905 65.125 ;
        RECT 9.095 64.955 9.995 65.125 ;
        RECT 10.285 64.955 11.185 65.125 ;
        RECT 11.475 64.955 12.375 65.125 ;
        RECT 12.665 64.955 13.565 65.125 ;
        RECT 13.855 64.955 14.755 65.125 ;
      LAYER mcon ;
        RECT 1.325 75.505 2.065 75.675 ;
        RECT 2.515 75.505 3.255 75.675 ;
        RECT 3.705 75.505 4.445 75.675 ;
        RECT 4.895 75.505 5.635 75.675 ;
        RECT 6.085 75.505 6.825 75.675 ;
        RECT 9.175 75.505 9.915 75.675 ;
        RECT 10.365 75.505 11.105 75.675 ;
        RECT 11.555 75.505 12.295 75.675 ;
        RECT 12.745 75.505 13.485 75.675 ;
        RECT 13.935 75.505 14.675 75.675 ;
        RECT 1.325 64.955 2.065 65.125 ;
        RECT 2.515 64.955 3.255 65.125 ;
        RECT 3.705 64.955 4.445 65.125 ;
        RECT 4.895 64.955 5.635 65.125 ;
        RECT 6.085 64.955 6.825 65.125 ;
        RECT 9.175 64.955 9.915 65.125 ;
        RECT 10.365 64.955 11.105 65.125 ;
        RECT 11.555 64.955 12.295 65.125 ;
        RECT 12.745 64.955 13.485 65.125 ;
        RECT 13.935 64.955 14.675 65.125 ;
      LAYER met1 ;
        RECT 2.470 75.980 14.735 75.985 ;
        RECT 0.110 75.475 14.735 75.980 ;
        RECT 0.110 75.470 2.470 75.475 ;
        RECT 0.110 65.155 0.620 75.470 ;
        RECT 0.110 64.645 14.735 65.155 ;
    END
  END in_hi
  PIN vss
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 15.700 102.560 18.480 105.050 ;
        RECT 15.700 95.050 23.535 102.560 ;
        RECT 14.145 82.470 24.025 95.050 ;
        RECT 0.105 64.025 15.895 76.605 ;
        RECT 24.335 71.405 34.215 95.065 ;
        RECT 34.275 71.405 73.555 95.065 ;
        RECT 1.875 59.700 14.265 63.800 ;
        RECT 16.825 60.550 23.475 68.130 ;
        RECT 14.145 46.780 24.025 59.360 ;
        RECT 15.700 39.270 23.535 46.780 ;
        RECT 24.335 46.765 34.215 70.425 ;
        RECT 34.275 46.765 73.555 70.425 ;
        RECT 15.700 36.780 18.480 39.270 ;
      LAYER li1 ;
        RECT 1.630 140.680 11.630 140.850 ;
        RECT 15.940 104.640 18.240 104.810 ;
        RECT 15.940 101.880 16.110 104.640 ;
        RECT 17.400 102.740 17.570 103.780 ;
        RECT 18.070 102.320 18.240 104.640 ;
        RECT 19.040 103.845 22.505 104.215 ;
        RECT 18.070 102.150 23.295 102.320 ;
        RECT 18.070 101.880 18.805 102.150 ;
        RECT 15.940 101.150 18.805 101.880 ;
        RECT 15.940 95.390 16.110 101.150 ;
        RECT 16.610 96.250 16.780 100.290 ;
        RECT 18.070 95.390 18.805 101.150 ;
        RECT 19.305 96.250 19.475 101.290 ;
        RECT 20.885 96.250 21.055 101.290 ;
        RECT 22.465 96.250 22.635 101.290 ;
        RECT 23.125 95.390 23.295 102.150 ;
        RECT 15.940 95.300 23.295 95.390 ;
        RECT 15.940 94.825 24.690 95.300 ;
        RECT 33.890 94.825 34.600 94.830 ;
        RECT 43.760 94.825 44.470 94.830 ;
        RECT 53.560 94.825 54.270 94.830 ;
        RECT 63.360 94.825 64.070 94.830 ;
        RECT 15.940 94.810 73.315 94.825 ;
        RECT 14.385 94.710 73.315 94.810 ;
        RECT 14.385 94.640 73.380 94.710 ;
        RECT 1.630 85.040 11.630 85.210 ;
        RECT 14.385 82.880 14.555 94.640 ;
        RECT 23.615 94.350 73.380 94.640 ;
        RECT 15.055 83.740 15.225 93.780 ;
        RECT 16.635 83.740 16.805 93.780 ;
        RECT 18.215 83.740 18.385 93.780 ;
        RECT 19.795 83.740 19.965 93.780 ;
        RECT 21.375 83.740 21.545 93.780 ;
        RECT 22.955 83.740 23.125 93.780 ;
        RECT 23.615 82.880 24.745 94.350 ;
        RECT 25.245 83.755 25.415 93.795 ;
        RECT 26.825 83.755 26.995 93.795 ;
        RECT 28.405 83.755 28.575 93.795 ;
        RECT 29.985 83.755 30.155 93.795 ;
        RECT 31.565 83.755 31.735 93.795 ;
        RECT 33.145 83.755 33.315 93.795 ;
        RECT 14.385 82.710 24.745 82.880 ;
        RECT 23.690 82.700 24.745 82.710 ;
        RECT 0.345 76.195 7.805 76.365 ;
        RECT 0.345 64.435 0.515 76.195 ;
        RECT 7.635 64.435 7.805 76.195 ;
        RECT 0.345 64.425 7.805 64.435 ;
        RECT 8.195 76.195 15.655 76.365 ;
        RECT 8.195 64.435 8.365 76.195 ;
        RECT 15.485 64.435 15.655 76.195 ;
        RECT 24.575 72.110 24.745 82.700 ;
        RECT 25.245 72.675 25.415 82.715 ;
        RECT 26.825 72.675 26.995 82.715 ;
        RECT 28.405 72.675 28.575 82.715 ;
        RECT 29.985 72.675 30.155 82.715 ;
        RECT 31.565 72.675 31.735 82.715 ;
        RECT 33.145 72.675 33.315 82.715 ;
        RECT 33.805 72.110 34.685 94.350 ;
        RECT 35.185 83.755 35.355 93.795 ;
        RECT 36.765 83.755 36.935 93.795 ;
        RECT 38.345 83.755 38.515 93.795 ;
        RECT 39.925 83.755 40.095 93.795 ;
        RECT 41.505 83.755 41.675 93.795 ;
        RECT 43.085 83.755 43.255 93.795 ;
        RECT 35.185 72.675 35.355 82.715 ;
        RECT 36.765 72.675 36.935 82.715 ;
        RECT 38.345 72.675 38.515 82.715 ;
        RECT 39.925 72.675 40.095 82.715 ;
        RECT 41.505 72.675 41.675 82.715 ;
        RECT 43.085 72.675 43.255 82.715 ;
        RECT 43.745 72.110 44.485 94.350 ;
        RECT 44.985 83.755 45.155 93.795 ;
        RECT 46.565 83.755 46.735 93.795 ;
        RECT 48.145 83.755 48.315 93.795 ;
        RECT 49.725 83.755 49.895 93.795 ;
        RECT 51.305 83.755 51.475 93.795 ;
        RECT 52.885 83.755 53.055 93.795 ;
        RECT 44.985 72.675 45.155 82.715 ;
        RECT 46.565 72.675 46.735 82.715 ;
        RECT 48.145 72.675 48.315 82.715 ;
        RECT 49.725 72.675 49.895 82.715 ;
        RECT 51.305 72.675 51.475 82.715 ;
        RECT 52.885 72.675 53.055 82.715 ;
        RECT 53.545 72.110 54.285 94.350 ;
        RECT 54.785 83.755 54.955 93.795 ;
        RECT 56.365 83.755 56.535 93.795 ;
        RECT 57.945 83.755 58.115 93.795 ;
        RECT 59.525 83.755 59.695 93.795 ;
        RECT 61.105 83.755 61.275 93.795 ;
        RECT 62.685 83.755 62.855 93.795 ;
        RECT 54.785 72.675 54.955 82.715 ;
        RECT 56.365 72.675 56.535 82.715 ;
        RECT 57.945 72.675 58.115 82.715 ;
        RECT 59.525 72.675 59.695 82.715 ;
        RECT 61.105 72.675 61.275 82.715 ;
        RECT 62.685 72.675 62.855 82.715 ;
        RECT 63.345 72.110 64.085 94.350 ;
        RECT 64.585 83.755 64.755 93.795 ;
        RECT 66.165 83.755 66.335 93.795 ;
        RECT 67.745 83.755 67.915 93.795 ;
        RECT 69.325 83.755 69.495 93.795 ;
        RECT 70.905 83.755 71.075 93.795 ;
        RECT 72.485 83.755 72.655 93.795 ;
        RECT 64.585 72.675 64.755 82.715 ;
        RECT 66.165 72.675 66.335 82.715 ;
        RECT 67.745 72.675 67.915 82.715 ;
        RECT 69.325 72.675 69.495 82.715 ;
        RECT 70.905 72.675 71.075 82.715 ;
        RECT 72.485 72.675 72.655 82.715 ;
        RECT 73.145 72.110 73.315 94.350 ;
        RECT 24.575 71.750 73.340 72.110 ;
        RECT 24.575 71.645 73.315 71.750 ;
        RECT 33.890 71.640 34.600 71.645 ;
        RECT 43.760 71.640 44.470 71.645 ;
        RECT 53.560 71.640 54.270 71.645 ;
        RECT 63.360 71.640 64.070 71.645 ;
        RECT 33.890 70.185 34.600 70.190 ;
        RECT 43.760 70.185 44.470 70.190 ;
        RECT 53.560 70.185 54.270 70.190 ;
        RECT 63.360 70.185 64.070 70.190 ;
        RECT 24.575 70.080 73.315 70.185 ;
        RECT 24.575 69.720 73.340 70.080 ;
        RECT 8.195 64.425 15.655 64.435 ;
        RECT 0.345 64.265 15.655 64.425 ;
        RECT 17.065 67.720 23.235 67.890 ;
        RECT 2.025 63.495 14.095 64.265 ;
        RECT 2.055 63.450 14.085 63.495 ;
        RECT 2.055 60.050 2.225 63.450 ;
        RECT 2.625 60.730 2.795 62.770 ;
        RECT 3.585 60.730 3.755 62.770 ;
        RECT 4.545 60.730 4.715 62.770 ;
        RECT 5.495 60.730 5.665 62.770 ;
        RECT 6.455 60.730 6.625 62.770 ;
        RECT 7.415 60.730 7.585 62.770 ;
        RECT 7.985 61.425 8.155 63.450 ;
        RECT 7.925 60.805 8.205 61.425 ;
        RECT 7.985 60.050 8.155 60.805 ;
        RECT 8.555 60.730 8.725 62.770 ;
        RECT 9.515 60.730 9.685 62.770 ;
        RECT 10.475 60.730 10.645 62.770 ;
        RECT 11.425 60.730 11.595 62.770 ;
        RECT 12.385 60.730 12.555 62.770 ;
        RECT 13.345 60.730 13.515 62.770 ;
        RECT 13.915 60.050 14.085 63.450 ;
        RECT 17.065 60.960 17.235 67.720 ;
        RECT 17.735 61.820 17.905 66.860 ;
        RECT 19.315 61.820 19.485 66.860 ;
        RECT 19.985 62.880 20.315 67.720 ;
        RECT 19.935 62.030 20.355 62.880 ;
        RECT 19.985 60.960 20.315 62.030 ;
        RECT 20.815 61.820 20.985 66.860 ;
        RECT 22.395 61.820 22.565 66.860 ;
        RECT 23.065 60.960 23.235 67.720 ;
        RECT 17.065 60.790 23.235 60.960 ;
        RECT 2.055 59.880 14.085 60.050 ;
        RECT 24.575 59.130 24.745 69.720 ;
        RECT 23.690 59.120 24.745 59.130 ;
        RECT 14.385 58.950 24.745 59.120 ;
        RECT 25.245 59.115 25.415 69.155 ;
        RECT 26.825 59.115 26.995 69.155 ;
        RECT 28.405 59.115 28.575 69.155 ;
        RECT 29.985 59.115 30.155 69.155 ;
        RECT 31.565 59.115 31.735 69.155 ;
        RECT 33.145 59.115 33.315 69.155 ;
        RECT 1.530 56.720 11.530 56.890 ;
        RECT 14.385 47.190 14.555 58.950 ;
        RECT 15.055 48.050 15.225 58.090 ;
        RECT 16.635 48.050 16.805 58.090 ;
        RECT 18.215 48.050 18.385 58.090 ;
        RECT 19.795 48.050 19.965 58.090 ;
        RECT 21.375 48.050 21.545 58.090 ;
        RECT 22.955 48.050 23.125 58.090 ;
        RECT 23.615 47.480 24.745 58.950 ;
        RECT 25.245 48.035 25.415 58.075 ;
        RECT 26.825 48.035 26.995 58.075 ;
        RECT 28.405 48.035 28.575 58.075 ;
        RECT 29.985 48.035 30.155 58.075 ;
        RECT 31.565 48.035 31.735 58.075 ;
        RECT 33.145 48.035 33.315 58.075 ;
        RECT 33.805 47.480 34.685 69.720 ;
        RECT 35.185 59.115 35.355 69.155 ;
        RECT 36.765 59.115 36.935 69.155 ;
        RECT 38.345 59.115 38.515 69.155 ;
        RECT 39.925 59.115 40.095 69.155 ;
        RECT 41.505 59.115 41.675 69.155 ;
        RECT 43.085 59.115 43.255 69.155 ;
        RECT 35.185 48.035 35.355 58.075 ;
        RECT 36.765 48.035 36.935 58.075 ;
        RECT 38.345 48.035 38.515 58.075 ;
        RECT 39.925 48.035 40.095 58.075 ;
        RECT 41.505 48.035 41.675 58.075 ;
        RECT 43.085 48.035 43.255 58.075 ;
        RECT 43.745 47.480 44.485 69.720 ;
        RECT 44.985 59.115 45.155 69.155 ;
        RECT 46.565 59.115 46.735 69.155 ;
        RECT 48.145 59.115 48.315 69.155 ;
        RECT 49.725 59.115 49.895 69.155 ;
        RECT 51.305 59.115 51.475 69.155 ;
        RECT 52.885 59.115 53.055 69.155 ;
        RECT 44.985 48.035 45.155 58.075 ;
        RECT 46.565 48.035 46.735 58.075 ;
        RECT 48.145 48.035 48.315 58.075 ;
        RECT 49.725 48.035 49.895 58.075 ;
        RECT 51.305 48.035 51.475 58.075 ;
        RECT 52.885 48.035 53.055 58.075 ;
        RECT 53.545 47.480 54.285 69.720 ;
        RECT 54.785 59.115 54.955 69.155 ;
        RECT 56.365 59.115 56.535 69.155 ;
        RECT 57.945 59.115 58.115 69.155 ;
        RECT 59.525 59.115 59.695 69.155 ;
        RECT 61.105 59.115 61.275 69.155 ;
        RECT 62.685 59.115 62.855 69.155 ;
        RECT 54.785 48.035 54.955 58.075 ;
        RECT 56.365 48.035 56.535 58.075 ;
        RECT 57.945 48.035 58.115 58.075 ;
        RECT 59.525 48.035 59.695 58.075 ;
        RECT 61.105 48.035 61.275 58.075 ;
        RECT 62.685 48.035 62.855 58.075 ;
        RECT 63.345 47.480 64.085 69.720 ;
        RECT 64.585 59.115 64.755 69.155 ;
        RECT 66.165 59.115 66.335 69.155 ;
        RECT 67.745 59.115 67.915 69.155 ;
        RECT 69.325 59.115 69.495 69.155 ;
        RECT 70.905 59.115 71.075 69.155 ;
        RECT 72.485 59.115 72.655 69.155 ;
        RECT 64.585 48.035 64.755 58.075 ;
        RECT 66.165 48.035 66.335 58.075 ;
        RECT 67.745 48.035 67.915 58.075 ;
        RECT 69.325 48.035 69.495 58.075 ;
        RECT 70.905 48.035 71.075 58.075 ;
        RECT 72.485 48.035 72.655 58.075 ;
        RECT 73.145 47.480 73.315 69.720 ;
        RECT 23.615 47.190 73.380 47.480 ;
        RECT 14.385 47.120 73.380 47.190 ;
        RECT 14.385 47.020 73.315 47.120 ;
        RECT 15.940 47.005 73.315 47.020 ;
        RECT 15.940 46.530 24.690 47.005 ;
        RECT 33.890 47.000 34.600 47.005 ;
        RECT 43.760 47.000 44.470 47.005 ;
        RECT 53.560 47.000 54.270 47.005 ;
        RECT 63.360 47.000 64.070 47.005 ;
        RECT 15.940 46.440 23.295 46.530 ;
        RECT 15.940 40.680 16.110 46.440 ;
        RECT 16.610 41.540 16.780 45.580 ;
        RECT 18.070 40.680 18.805 46.440 ;
        RECT 15.940 39.950 18.805 40.680 ;
        RECT 19.305 40.540 19.475 45.580 ;
        RECT 20.885 40.540 21.055 45.580 ;
        RECT 22.465 40.540 22.635 45.580 ;
        RECT 15.940 37.190 16.110 39.950 ;
        RECT 18.070 39.680 18.805 39.950 ;
        RECT 23.125 39.680 23.295 46.440 ;
        RECT 18.070 39.510 23.295 39.680 ;
        RECT 17.400 38.050 17.570 39.090 ;
        RECT 18.070 37.190 18.240 39.510 ;
        RECT 19.040 37.615 22.505 37.985 ;
        RECT 15.940 37.020 18.240 37.190 ;
        RECT 1.530 1.080 11.530 1.250 ;
      LAYER mcon ;
        RECT 1.710 140.680 11.550 140.850 ;
        RECT 17.400 102.820 17.570 103.700 ;
        RECT 19.070 103.875 19.380 104.185 ;
        RECT 22.135 103.845 22.505 104.215 ;
        RECT 16.610 96.330 16.780 100.210 ;
        RECT 19.305 96.330 19.475 101.210 ;
        RECT 20.885 96.330 21.055 101.210 ;
        RECT 22.465 96.330 22.635 101.210 ;
        RECT 1.710 85.040 11.550 85.210 ;
        RECT 15.055 83.820 15.225 93.700 ;
        RECT 16.635 83.820 16.805 93.700 ;
        RECT 18.215 83.820 18.385 93.700 ;
        RECT 19.795 83.820 19.965 93.700 ;
        RECT 21.375 83.820 21.545 93.700 ;
        RECT 22.955 83.820 23.125 93.700 ;
        RECT 25.245 83.835 25.415 93.715 ;
        RECT 26.825 83.835 26.995 93.715 ;
        RECT 28.405 83.835 28.575 93.715 ;
        RECT 29.985 83.835 30.155 93.715 ;
        RECT 31.565 83.835 31.735 93.715 ;
        RECT 33.145 83.835 33.315 93.715 ;
        RECT 25.245 72.755 25.415 82.635 ;
        RECT 26.825 72.755 26.995 82.635 ;
        RECT 28.405 72.755 28.575 82.635 ;
        RECT 29.985 72.755 30.155 82.635 ;
        RECT 31.565 72.755 31.735 82.635 ;
        RECT 33.145 72.755 33.315 82.635 ;
        RECT 35.185 83.835 35.355 93.715 ;
        RECT 36.765 83.835 36.935 93.715 ;
        RECT 38.345 83.835 38.515 93.715 ;
        RECT 39.925 83.835 40.095 93.715 ;
        RECT 41.505 83.835 41.675 93.715 ;
        RECT 43.085 83.835 43.255 93.715 ;
        RECT 43.770 84.970 44.460 87.390 ;
        RECT 33.900 73.840 34.590 76.260 ;
        RECT 35.185 72.755 35.355 82.635 ;
        RECT 36.765 72.755 36.935 82.635 ;
        RECT 38.345 72.755 38.515 82.635 ;
        RECT 39.925 72.755 40.095 82.635 ;
        RECT 41.505 72.755 41.675 82.635 ;
        RECT 43.085 72.755 43.255 82.635 ;
        RECT 44.985 83.835 45.155 93.715 ;
        RECT 46.565 83.835 46.735 93.715 ;
        RECT 48.145 83.835 48.315 93.715 ;
        RECT 49.725 83.835 49.895 93.715 ;
        RECT 51.305 83.835 51.475 93.715 ;
        RECT 52.885 83.835 53.055 93.715 ;
        RECT 44.985 72.755 45.155 82.635 ;
        RECT 46.565 72.755 46.735 82.635 ;
        RECT 48.145 72.755 48.315 82.635 ;
        RECT 49.725 72.755 49.895 82.635 ;
        RECT 51.305 72.755 51.475 82.635 ;
        RECT 52.885 72.755 53.055 82.635 ;
        RECT 54.785 83.835 54.955 93.715 ;
        RECT 56.365 83.835 56.535 93.715 ;
        RECT 57.945 83.835 58.115 93.715 ;
        RECT 59.525 83.835 59.695 93.715 ;
        RECT 61.105 83.835 61.275 93.715 ;
        RECT 62.685 83.835 62.855 93.715 ;
        RECT 63.350 84.970 64.040 87.390 ;
        RECT 53.570 73.850 54.260 76.270 ;
        RECT 54.785 72.755 54.955 82.635 ;
        RECT 56.365 72.755 56.535 82.635 ;
        RECT 57.945 72.755 58.115 82.635 ;
        RECT 59.525 72.755 59.695 82.635 ;
        RECT 61.105 72.755 61.275 82.635 ;
        RECT 62.685 72.755 62.855 82.635 ;
        RECT 64.585 83.835 64.755 93.715 ;
        RECT 66.165 83.835 66.335 93.715 ;
        RECT 67.745 83.835 67.915 93.715 ;
        RECT 69.325 83.835 69.495 93.715 ;
        RECT 70.905 83.835 71.075 93.715 ;
        RECT 72.485 83.835 72.655 93.715 ;
        RECT 64.585 72.755 64.755 82.635 ;
        RECT 66.165 72.755 66.335 82.635 ;
        RECT 67.745 72.755 67.915 82.635 ;
        RECT 69.325 72.755 69.495 82.635 ;
        RECT 70.905 72.755 71.075 82.635 ;
        RECT 72.485 72.755 72.655 82.635 ;
        RECT 2.625 60.810 2.795 62.690 ;
        RECT 3.585 60.810 3.755 62.690 ;
        RECT 4.545 60.810 4.715 62.690 ;
        RECT 5.495 60.810 5.665 62.690 ;
        RECT 6.455 60.810 6.625 62.690 ;
        RECT 7.415 60.810 7.585 62.690 ;
        RECT 7.925 60.805 8.205 61.425 ;
        RECT 8.555 60.810 8.725 62.690 ;
        RECT 9.515 60.810 9.685 62.690 ;
        RECT 10.475 60.810 10.645 62.690 ;
        RECT 11.425 60.810 11.595 62.690 ;
        RECT 12.385 60.810 12.555 62.690 ;
        RECT 13.345 60.810 13.515 62.690 ;
        RECT 17.735 61.900 17.905 66.780 ;
        RECT 19.315 61.900 19.485 66.780 ;
        RECT 19.935 62.030 20.355 62.880 ;
        RECT 20.815 61.900 20.985 66.780 ;
        RECT 22.395 61.900 22.565 66.780 ;
        RECT 25.245 59.195 25.415 69.075 ;
        RECT 26.825 59.195 26.995 69.075 ;
        RECT 28.405 59.195 28.575 69.075 ;
        RECT 29.985 59.195 30.155 69.075 ;
        RECT 31.565 59.195 31.735 69.075 ;
        RECT 33.145 59.195 33.315 69.075 ;
        RECT 33.900 65.570 34.590 67.990 ;
        RECT 1.610 56.720 11.450 56.890 ;
        RECT 15.055 48.130 15.225 58.010 ;
        RECT 16.635 48.130 16.805 58.010 ;
        RECT 18.215 48.130 18.385 58.010 ;
        RECT 19.795 48.130 19.965 58.010 ;
        RECT 21.375 48.130 21.545 58.010 ;
        RECT 22.955 48.130 23.125 58.010 ;
        RECT 25.245 48.115 25.415 57.995 ;
        RECT 26.825 48.115 26.995 57.995 ;
        RECT 28.405 48.115 28.575 57.995 ;
        RECT 29.985 48.115 30.155 57.995 ;
        RECT 31.565 48.115 31.735 57.995 ;
        RECT 33.145 48.115 33.315 57.995 ;
        RECT 35.185 59.195 35.355 69.075 ;
        RECT 36.765 59.195 36.935 69.075 ;
        RECT 38.345 59.195 38.515 69.075 ;
        RECT 39.925 59.195 40.095 69.075 ;
        RECT 41.505 59.195 41.675 69.075 ;
        RECT 43.085 59.195 43.255 69.075 ;
        RECT 35.185 48.115 35.355 57.995 ;
        RECT 36.765 48.115 36.935 57.995 ;
        RECT 38.345 48.115 38.515 57.995 ;
        RECT 39.925 48.115 40.095 57.995 ;
        RECT 41.505 48.115 41.675 57.995 ;
        RECT 43.085 48.115 43.255 57.995 ;
        RECT 44.985 59.195 45.155 69.075 ;
        RECT 46.565 59.195 46.735 69.075 ;
        RECT 48.145 59.195 48.315 69.075 ;
        RECT 49.725 59.195 49.895 69.075 ;
        RECT 51.305 59.195 51.475 69.075 ;
        RECT 52.885 59.195 53.055 69.075 ;
        RECT 53.570 65.560 54.260 67.980 ;
        RECT 43.770 54.440 44.460 56.860 ;
        RECT 44.985 48.115 45.155 57.995 ;
        RECT 46.565 48.115 46.735 57.995 ;
        RECT 48.145 48.115 48.315 57.995 ;
        RECT 49.725 48.115 49.895 57.995 ;
        RECT 51.305 48.115 51.475 57.995 ;
        RECT 52.885 48.115 53.055 57.995 ;
        RECT 54.785 59.195 54.955 69.075 ;
        RECT 56.365 59.195 56.535 69.075 ;
        RECT 57.945 59.195 58.115 69.075 ;
        RECT 59.525 59.195 59.695 69.075 ;
        RECT 61.105 59.195 61.275 69.075 ;
        RECT 62.685 59.195 62.855 69.075 ;
        RECT 54.785 48.115 54.955 57.995 ;
        RECT 56.365 48.115 56.535 57.995 ;
        RECT 57.945 48.115 58.115 57.995 ;
        RECT 59.525 48.115 59.695 57.995 ;
        RECT 61.105 48.115 61.275 57.995 ;
        RECT 62.685 48.115 62.855 57.995 ;
        RECT 64.585 59.195 64.755 69.075 ;
        RECT 66.165 59.195 66.335 69.075 ;
        RECT 67.745 59.195 67.915 69.075 ;
        RECT 69.325 59.195 69.495 69.075 ;
        RECT 70.905 59.195 71.075 69.075 ;
        RECT 72.485 59.195 72.655 69.075 ;
        RECT 63.350 54.440 64.040 56.860 ;
        RECT 64.585 48.115 64.755 57.995 ;
        RECT 66.165 48.115 66.335 57.995 ;
        RECT 67.745 48.115 67.915 57.995 ;
        RECT 69.325 48.115 69.495 57.995 ;
        RECT 70.905 48.115 71.075 57.995 ;
        RECT 72.485 48.115 72.655 57.995 ;
        RECT 16.610 41.620 16.780 45.500 ;
        RECT 19.305 40.620 19.475 45.500 ;
        RECT 20.885 40.620 21.055 45.500 ;
        RECT 22.465 40.620 22.635 45.500 ;
        RECT 17.400 38.130 17.570 39.010 ;
        RECT 19.070 37.645 19.380 37.955 ;
        RECT 22.135 37.615 22.505 37.985 ;
        RECT 1.610 1.080 11.450 1.250 ;
      LAYER met1 ;
        RECT 1.650 140.650 11.610 140.880 ;
        RECT 17.370 103.740 17.600 103.760 ;
        RECT 18.820 103.740 19.480 104.270 ;
        RECT 17.370 103.370 19.480 103.740 ;
        RECT 17.370 102.760 17.600 103.370 ;
        RECT 21.940 103.030 22.720 104.390 ;
        RECT 16.580 97.290 16.810 100.270 ;
        RECT 16.440 96.620 16.890 97.290 ;
        RECT 19.275 97.280 19.505 101.270 ;
        RECT 20.855 97.290 21.085 101.270 ;
        RECT 19.190 96.630 19.590 97.280 ;
        RECT 20.790 96.640 21.190 97.290 ;
        RECT 22.435 97.260 22.665 101.270 ;
        RECT 16.580 96.270 16.810 96.620 ;
        RECT 19.275 96.270 19.505 96.630 ;
        RECT 20.855 96.270 21.085 96.640 ;
        RECT 22.340 96.610 22.740 97.260 ;
        RECT 22.435 96.270 22.665 96.610 ;
        RECT 1.570 84.640 11.660 85.240 ;
        RECT 15.025 84.990 15.255 93.760 ;
        RECT 14.930 84.340 15.330 84.990 ;
        RECT 16.605 84.980 16.835 93.760 ;
        RECT 18.185 84.980 18.415 93.760 ;
        RECT 19.765 84.980 19.995 93.760 ;
        RECT 21.345 84.980 21.575 93.760 ;
        RECT 22.925 84.980 23.155 93.760 ;
        RECT 25.215 88.370 25.445 93.775 ;
        RECT 26.795 88.370 27.025 93.775 ;
        RECT 15.025 83.760 15.255 84.340 ;
        RECT 16.510 84.330 16.910 84.980 ;
        RECT 18.100 84.330 18.500 84.980 ;
        RECT 19.680 84.330 20.080 84.980 ;
        RECT 21.260 84.330 21.660 84.980 ;
        RECT 22.850 84.330 23.250 84.980 ;
        RECT 16.605 83.760 16.835 84.330 ;
        RECT 18.185 83.760 18.415 84.330 ;
        RECT 19.765 83.760 19.995 84.330 ;
        RECT 21.345 83.760 21.575 84.330 ;
        RECT 22.925 83.760 23.155 84.330 ;
        RECT 24.950 84.020 25.680 88.370 ;
        RECT 26.540 84.020 27.270 88.370 ;
        RECT 28.375 88.360 28.605 93.775 ;
        RECT 29.955 88.360 30.185 93.775 ;
        RECT 31.535 88.360 31.765 93.775 ;
        RECT 33.115 88.360 33.345 93.775 ;
        RECT 35.155 88.370 35.385 93.775 ;
        RECT 36.735 88.370 36.965 93.775 ;
        RECT 25.215 83.775 25.445 84.020 ;
        RECT 26.795 83.775 27.025 84.020 ;
        RECT 28.110 84.010 28.840 88.360 ;
        RECT 29.690 84.010 30.420 88.360 ;
        RECT 31.280 84.010 32.010 88.360 ;
        RECT 32.850 84.010 33.580 88.360 ;
        RECT 34.880 84.020 35.610 88.370 ;
        RECT 36.470 84.020 37.200 88.370 ;
        RECT 38.315 88.360 38.545 93.775 ;
        RECT 39.895 88.360 40.125 93.775 ;
        RECT 41.475 88.360 41.705 93.775 ;
        RECT 43.055 88.360 43.285 93.775 ;
        RECT 44.955 88.370 45.185 93.775 ;
        RECT 46.535 88.370 46.765 93.775 ;
        RECT 28.375 83.775 28.605 84.010 ;
        RECT 29.955 83.775 30.185 84.010 ;
        RECT 31.535 83.775 31.765 84.010 ;
        RECT 33.115 83.775 33.345 84.010 ;
        RECT 35.155 83.775 35.385 84.020 ;
        RECT 36.735 83.775 36.965 84.020 ;
        RECT 38.040 84.010 38.770 88.360 ;
        RECT 39.620 84.010 40.350 88.360 ;
        RECT 41.210 84.010 41.940 88.360 ;
        RECT 42.780 84.010 43.510 88.360 ;
        RECT 43.740 87.390 44.490 87.450 ;
        RECT 43.720 84.970 44.510 87.390 ;
        RECT 43.740 84.910 44.490 84.970 ;
        RECT 44.690 84.020 45.420 88.370 ;
        RECT 46.280 84.020 47.010 88.370 ;
        RECT 48.115 88.360 48.345 93.775 ;
        RECT 49.695 88.360 49.925 93.775 ;
        RECT 51.275 88.360 51.505 93.775 ;
        RECT 52.855 88.360 53.085 93.775 ;
        RECT 38.315 83.775 38.545 84.010 ;
        RECT 39.895 83.775 40.125 84.010 ;
        RECT 41.475 83.775 41.705 84.010 ;
        RECT 43.055 83.775 43.285 84.010 ;
        RECT 44.955 83.775 45.185 84.020 ;
        RECT 46.535 83.775 46.765 84.020 ;
        RECT 47.850 84.010 48.580 88.360 ;
        RECT 49.430 84.010 50.160 88.360 ;
        RECT 51.020 84.010 51.750 88.360 ;
        RECT 52.590 84.010 53.320 88.360 ;
        RECT 54.755 88.340 54.985 93.775 ;
        RECT 56.335 88.340 56.565 93.775 ;
        RECT 48.115 83.775 48.345 84.010 ;
        RECT 49.695 83.775 49.925 84.010 ;
        RECT 51.275 83.775 51.505 84.010 ;
        RECT 52.855 83.775 53.085 84.010 ;
        RECT 54.500 83.990 55.230 88.340 ;
        RECT 56.090 83.990 56.820 88.340 ;
        RECT 57.915 88.330 58.145 93.775 ;
        RECT 59.495 88.330 59.725 93.775 ;
        RECT 61.075 88.330 61.305 93.775 ;
        RECT 62.655 88.330 62.885 93.775 ;
        RECT 64.555 88.340 64.785 93.775 ;
        RECT 66.135 88.340 66.365 93.775 ;
        RECT 54.755 83.775 54.985 83.990 ;
        RECT 56.335 83.775 56.565 83.990 ;
        RECT 57.660 83.980 58.390 88.330 ;
        RECT 59.240 83.980 59.970 88.330 ;
        RECT 60.830 83.980 61.560 88.330 ;
        RECT 62.400 83.980 63.130 88.330 ;
        RECT 63.320 87.390 64.070 87.450 ;
        RECT 63.300 84.970 64.090 87.390 ;
        RECT 63.320 84.910 64.070 84.970 ;
        RECT 64.290 83.990 65.020 88.340 ;
        RECT 65.880 83.990 66.610 88.340 ;
        RECT 67.715 88.330 67.945 93.775 ;
        RECT 69.295 88.330 69.525 93.775 ;
        RECT 70.875 88.330 71.105 93.775 ;
        RECT 72.455 88.330 72.685 93.775 ;
        RECT 57.915 83.775 58.145 83.980 ;
        RECT 59.495 83.775 59.725 83.980 ;
        RECT 61.075 83.775 61.305 83.980 ;
        RECT 62.655 83.775 62.885 83.980 ;
        RECT 64.555 83.775 64.785 83.990 ;
        RECT 66.135 83.775 66.365 83.990 ;
        RECT 67.450 83.980 68.180 88.330 ;
        RECT 69.030 83.980 69.760 88.330 ;
        RECT 70.620 83.980 71.350 88.330 ;
        RECT 72.190 83.980 72.920 88.330 ;
        RECT 67.715 83.775 67.945 83.980 ;
        RECT 69.295 83.775 69.525 83.980 ;
        RECT 70.875 83.775 71.105 83.980 ;
        RECT 72.455 83.775 72.685 83.980 ;
        RECT 25.215 77.320 25.445 82.695 ;
        RECT 26.795 77.320 27.025 82.695 ;
        RECT 24.960 72.970 25.690 77.320 ;
        RECT 26.550 72.970 27.280 77.320 ;
        RECT 28.375 77.310 28.605 82.695 ;
        RECT 29.955 77.310 30.185 82.695 ;
        RECT 31.535 77.310 31.765 82.695 ;
        RECT 33.115 77.310 33.345 82.695 ;
        RECT 35.155 77.320 35.385 82.695 ;
        RECT 36.735 77.320 36.965 82.695 ;
        RECT 25.215 72.695 25.445 72.970 ;
        RECT 26.795 72.695 27.025 72.970 ;
        RECT 28.120 72.960 28.850 77.310 ;
        RECT 29.700 72.960 30.430 77.310 ;
        RECT 31.290 72.960 32.020 77.310 ;
        RECT 32.860 72.960 33.590 77.310 ;
        RECT 33.870 76.260 34.620 76.320 ;
        RECT 33.850 73.840 34.640 76.260 ;
        RECT 33.870 73.780 34.620 73.840 ;
        RECT 34.890 72.970 35.620 77.320 ;
        RECT 36.480 72.970 37.210 77.320 ;
        RECT 38.315 77.310 38.545 82.695 ;
        RECT 39.895 77.310 40.125 82.695 ;
        RECT 41.475 77.310 41.705 82.695 ;
        RECT 43.055 77.310 43.285 82.695 ;
        RECT 44.955 77.320 45.185 82.695 ;
        RECT 46.535 77.320 46.765 82.695 ;
        RECT 28.375 72.695 28.605 72.960 ;
        RECT 29.955 72.695 30.185 72.960 ;
        RECT 31.535 72.695 31.765 72.960 ;
        RECT 33.115 72.695 33.345 72.960 ;
        RECT 35.155 72.695 35.385 72.970 ;
        RECT 36.735 72.695 36.965 72.970 ;
        RECT 38.050 72.960 38.780 77.310 ;
        RECT 39.630 72.960 40.360 77.310 ;
        RECT 41.220 72.960 41.950 77.310 ;
        RECT 42.790 72.960 43.520 77.310 ;
        RECT 44.700 72.970 45.430 77.320 ;
        RECT 46.290 72.970 47.020 77.320 ;
        RECT 48.115 77.310 48.345 82.695 ;
        RECT 49.695 77.310 49.925 82.695 ;
        RECT 51.275 77.310 51.505 82.695 ;
        RECT 52.855 77.310 53.085 82.695 ;
        RECT 38.315 72.695 38.545 72.960 ;
        RECT 39.895 72.695 40.125 72.960 ;
        RECT 41.475 72.695 41.705 72.960 ;
        RECT 43.055 72.695 43.285 72.960 ;
        RECT 44.955 72.695 45.185 72.970 ;
        RECT 46.535 72.695 46.765 72.970 ;
        RECT 47.860 72.960 48.590 77.310 ;
        RECT 49.440 72.960 50.170 77.310 ;
        RECT 51.030 72.960 51.760 77.310 ;
        RECT 52.600 72.960 53.330 77.310 ;
        RECT 54.755 77.290 54.985 82.695 ;
        RECT 56.335 77.290 56.565 82.695 ;
        RECT 53.540 76.270 54.290 76.330 ;
        RECT 53.520 73.850 54.310 76.270 ;
        RECT 53.540 73.790 54.290 73.850 ;
        RECT 48.115 72.695 48.345 72.960 ;
        RECT 49.695 72.695 49.925 72.960 ;
        RECT 51.275 72.695 51.505 72.960 ;
        RECT 52.855 72.695 53.085 72.960 ;
        RECT 54.510 72.940 55.240 77.290 ;
        RECT 56.100 72.940 56.830 77.290 ;
        RECT 57.915 77.280 58.145 82.695 ;
        RECT 59.495 77.280 59.725 82.695 ;
        RECT 61.075 77.280 61.305 82.695 ;
        RECT 62.655 77.280 62.885 82.695 ;
        RECT 64.555 77.290 64.785 82.695 ;
        RECT 66.135 77.290 66.365 82.695 ;
        RECT 54.755 72.695 54.985 72.940 ;
        RECT 56.335 72.695 56.565 72.940 ;
        RECT 57.670 72.930 58.400 77.280 ;
        RECT 59.250 72.930 59.980 77.280 ;
        RECT 60.840 72.930 61.570 77.280 ;
        RECT 62.410 72.930 63.140 77.280 ;
        RECT 64.300 72.940 65.030 77.290 ;
        RECT 65.890 72.940 66.620 77.290 ;
        RECT 67.715 77.280 67.945 82.695 ;
        RECT 69.295 77.280 69.525 82.695 ;
        RECT 70.875 77.280 71.105 82.695 ;
        RECT 72.455 77.280 72.685 82.695 ;
        RECT 57.915 72.695 58.145 72.930 ;
        RECT 59.495 72.695 59.725 72.930 ;
        RECT 61.075 72.695 61.305 72.930 ;
        RECT 62.655 72.695 62.885 72.930 ;
        RECT 64.555 72.695 64.785 72.940 ;
        RECT 66.135 72.695 66.365 72.940 ;
        RECT 67.460 72.930 68.190 77.280 ;
        RECT 69.040 72.930 69.770 77.280 ;
        RECT 70.630 72.930 71.360 77.280 ;
        RECT 72.200 72.930 72.930 77.280 ;
        RECT 67.715 72.695 67.945 72.930 ;
        RECT 69.295 72.695 69.525 72.930 ;
        RECT 70.875 72.695 71.105 72.930 ;
        RECT 72.455 72.695 72.685 72.930 ;
        RECT 25.215 68.860 25.445 69.135 ;
        RECT 26.795 68.860 27.025 69.135 ;
        RECT 28.375 68.870 28.605 69.135 ;
        RECT 29.955 68.870 30.185 69.135 ;
        RECT 31.535 68.870 31.765 69.135 ;
        RECT 33.115 68.870 33.345 69.135 ;
        RECT 17.705 62.880 17.935 66.840 ;
        RECT 19.285 62.880 19.515 66.840 ;
        RECT 19.905 62.880 20.385 62.940 ;
        RECT 20.785 62.880 21.015 66.840 ;
        RECT 22.365 62.880 22.595 66.840 ;
        RECT 24.960 64.510 25.690 68.860 ;
        RECT 26.550 64.510 27.280 68.860 ;
        RECT 28.120 64.520 28.850 68.870 ;
        RECT 29.700 64.520 30.430 68.870 ;
        RECT 31.290 64.520 32.020 68.870 ;
        RECT 32.860 64.520 33.590 68.870 ;
        RECT 35.155 68.860 35.385 69.135 ;
        RECT 36.735 68.860 36.965 69.135 ;
        RECT 38.315 68.870 38.545 69.135 ;
        RECT 39.895 68.870 40.125 69.135 ;
        RECT 41.475 68.870 41.705 69.135 ;
        RECT 43.055 68.870 43.285 69.135 ;
        RECT 33.870 67.990 34.620 68.050 ;
        RECT 33.850 65.570 34.640 67.990 ;
        RECT 33.870 65.510 34.620 65.570 ;
        RECT 2.595 61.425 2.825 62.750 ;
        RECT 3.555 61.425 3.785 62.750 ;
        RECT 4.515 61.425 4.745 62.750 ;
        RECT 5.465 61.425 5.695 62.750 ;
        RECT 6.425 61.425 6.655 62.750 ;
        RECT 7.385 61.425 7.615 62.750 ;
        RECT 7.895 61.425 8.235 61.485 ;
        RECT 8.525 61.425 8.755 62.750 ;
        RECT 9.485 61.425 9.715 62.750 ;
        RECT 10.445 61.425 10.675 62.750 ;
        RECT 11.395 61.425 11.625 62.750 ;
        RECT 12.355 61.425 12.585 62.750 ;
        RECT 13.315 61.425 13.545 62.750 ;
        RECT 17.645 62.030 18.005 62.880 ;
        RECT 19.225 62.030 19.585 62.880 ;
        RECT 19.885 62.030 20.405 62.880 ;
        RECT 20.725 62.030 21.085 62.880 ;
        RECT 22.295 62.030 22.655 62.880 ;
        RECT 17.705 61.840 17.935 62.030 ;
        RECT 19.285 61.840 19.515 62.030 ;
        RECT 19.905 61.970 20.385 62.030 ;
        RECT 20.785 61.840 21.015 62.030 ;
        RECT 22.365 61.840 22.595 62.030 ;
        RECT 2.515 60.805 2.875 61.425 ;
        RECT 3.475 60.805 3.835 61.425 ;
        RECT 4.435 60.805 4.795 61.425 ;
        RECT 5.395 60.805 5.755 61.425 ;
        RECT 6.355 60.805 6.715 61.425 ;
        RECT 7.315 60.805 7.675 61.425 ;
        RECT 7.875 60.805 8.255 61.425 ;
        RECT 8.455 60.805 8.815 61.425 ;
        RECT 9.415 60.805 9.775 61.425 ;
        RECT 10.375 60.805 10.735 61.425 ;
        RECT 11.335 60.805 11.695 61.425 ;
        RECT 12.295 60.805 12.655 61.425 ;
        RECT 13.255 60.805 13.615 61.425 ;
        RECT 2.595 60.750 2.825 60.805 ;
        RECT 3.555 60.750 3.785 60.805 ;
        RECT 4.515 60.750 4.745 60.805 ;
        RECT 5.465 60.750 5.695 60.805 ;
        RECT 6.425 60.750 6.655 60.805 ;
        RECT 7.385 60.750 7.615 60.805 ;
        RECT 7.895 60.745 8.235 60.805 ;
        RECT 8.525 60.750 8.755 60.805 ;
        RECT 9.485 60.750 9.715 60.805 ;
        RECT 10.445 60.750 10.675 60.805 ;
        RECT 11.395 60.750 11.625 60.805 ;
        RECT 12.355 60.750 12.585 60.805 ;
        RECT 13.315 60.750 13.545 60.805 ;
        RECT 25.215 59.135 25.445 64.510 ;
        RECT 26.795 59.135 27.025 64.510 ;
        RECT 28.375 59.135 28.605 64.520 ;
        RECT 29.955 59.135 30.185 64.520 ;
        RECT 31.535 59.135 31.765 64.520 ;
        RECT 33.115 59.135 33.345 64.520 ;
        RECT 34.890 64.510 35.620 68.860 ;
        RECT 36.480 64.510 37.210 68.860 ;
        RECT 38.050 64.520 38.780 68.870 ;
        RECT 39.630 64.520 40.360 68.870 ;
        RECT 41.220 64.520 41.950 68.870 ;
        RECT 42.790 64.520 43.520 68.870 ;
        RECT 44.955 68.860 45.185 69.135 ;
        RECT 46.535 68.860 46.765 69.135 ;
        RECT 48.115 68.870 48.345 69.135 ;
        RECT 49.695 68.870 49.925 69.135 ;
        RECT 51.275 68.870 51.505 69.135 ;
        RECT 52.855 68.870 53.085 69.135 ;
        RECT 54.755 68.890 54.985 69.135 ;
        RECT 56.335 68.890 56.565 69.135 ;
        RECT 57.915 68.900 58.145 69.135 ;
        RECT 59.495 68.900 59.725 69.135 ;
        RECT 61.075 68.900 61.305 69.135 ;
        RECT 62.655 68.900 62.885 69.135 ;
        RECT 35.155 59.135 35.385 64.510 ;
        RECT 36.735 59.135 36.965 64.510 ;
        RECT 38.315 59.135 38.545 64.520 ;
        RECT 39.895 59.135 40.125 64.520 ;
        RECT 41.475 59.135 41.705 64.520 ;
        RECT 43.055 59.135 43.285 64.520 ;
        RECT 44.700 64.510 45.430 68.860 ;
        RECT 46.290 64.510 47.020 68.860 ;
        RECT 47.860 64.520 48.590 68.870 ;
        RECT 49.440 64.520 50.170 68.870 ;
        RECT 51.030 64.520 51.760 68.870 ;
        RECT 52.600 64.520 53.330 68.870 ;
        RECT 53.540 67.980 54.290 68.040 ;
        RECT 53.520 65.560 54.310 67.980 ;
        RECT 53.540 65.500 54.290 65.560 ;
        RECT 54.510 64.540 55.240 68.890 ;
        RECT 56.100 64.540 56.830 68.890 ;
        RECT 57.670 64.550 58.400 68.900 ;
        RECT 59.250 64.550 59.980 68.900 ;
        RECT 60.840 64.550 61.570 68.900 ;
        RECT 62.410 64.550 63.140 68.900 ;
        RECT 64.555 68.890 64.785 69.135 ;
        RECT 66.135 68.890 66.365 69.135 ;
        RECT 67.715 68.900 67.945 69.135 ;
        RECT 69.295 68.900 69.525 69.135 ;
        RECT 70.875 68.900 71.105 69.135 ;
        RECT 72.455 68.900 72.685 69.135 ;
        RECT 44.955 59.135 45.185 64.510 ;
        RECT 46.535 59.135 46.765 64.510 ;
        RECT 48.115 59.135 48.345 64.520 ;
        RECT 49.695 59.135 49.925 64.520 ;
        RECT 51.275 59.135 51.505 64.520 ;
        RECT 52.855 59.135 53.085 64.520 ;
        RECT 54.755 59.135 54.985 64.540 ;
        RECT 56.335 59.135 56.565 64.540 ;
        RECT 57.915 59.135 58.145 64.550 ;
        RECT 59.495 59.135 59.725 64.550 ;
        RECT 61.075 59.135 61.305 64.550 ;
        RECT 62.655 59.135 62.885 64.550 ;
        RECT 64.300 64.540 65.030 68.890 ;
        RECT 65.890 64.540 66.620 68.890 ;
        RECT 67.460 64.550 68.190 68.900 ;
        RECT 69.040 64.550 69.770 68.900 ;
        RECT 70.630 64.550 71.360 68.900 ;
        RECT 72.200 64.550 72.930 68.900 ;
        RECT 64.555 59.135 64.785 64.540 ;
        RECT 66.135 59.135 66.365 64.540 ;
        RECT 67.715 59.135 67.945 64.550 ;
        RECT 69.295 59.135 69.525 64.550 ;
        RECT 70.875 59.135 71.105 64.550 ;
        RECT 72.455 59.135 72.685 64.550 ;
        RECT 15.025 57.490 15.255 58.070 ;
        RECT 16.605 57.500 16.835 58.070 ;
        RECT 18.185 57.500 18.415 58.070 ;
        RECT 19.765 57.500 19.995 58.070 ;
        RECT 21.345 57.500 21.575 58.070 ;
        RECT 22.925 57.500 23.155 58.070 ;
        RECT 25.215 57.810 25.445 58.055 ;
        RECT 26.795 57.810 27.025 58.055 ;
        RECT 28.375 57.820 28.605 58.055 ;
        RECT 29.955 57.820 30.185 58.055 ;
        RECT 31.535 57.820 31.765 58.055 ;
        RECT 33.115 57.820 33.345 58.055 ;
        RECT 1.480 56.730 11.580 57.200 ;
        RECT 14.930 56.840 15.330 57.490 ;
        RECT 16.510 56.850 16.910 57.500 ;
        RECT 18.100 56.850 18.500 57.500 ;
        RECT 19.680 56.850 20.080 57.500 ;
        RECT 21.260 56.850 21.660 57.500 ;
        RECT 22.850 56.850 23.250 57.500 ;
        RECT 1.550 56.690 11.510 56.730 ;
        RECT 15.025 48.070 15.255 56.840 ;
        RECT 16.605 48.070 16.835 56.850 ;
        RECT 18.185 48.070 18.415 56.850 ;
        RECT 19.765 48.070 19.995 56.850 ;
        RECT 21.345 48.070 21.575 56.850 ;
        RECT 22.925 48.070 23.155 56.850 ;
        RECT 24.950 53.460 25.680 57.810 ;
        RECT 26.540 53.460 27.270 57.810 ;
        RECT 28.110 53.470 28.840 57.820 ;
        RECT 29.690 53.470 30.420 57.820 ;
        RECT 31.280 53.470 32.010 57.820 ;
        RECT 32.850 53.470 33.580 57.820 ;
        RECT 35.155 57.810 35.385 58.055 ;
        RECT 36.735 57.810 36.965 58.055 ;
        RECT 38.315 57.820 38.545 58.055 ;
        RECT 39.895 57.820 40.125 58.055 ;
        RECT 41.475 57.820 41.705 58.055 ;
        RECT 43.055 57.820 43.285 58.055 ;
        RECT 25.215 48.055 25.445 53.460 ;
        RECT 26.795 48.055 27.025 53.460 ;
        RECT 28.375 48.055 28.605 53.470 ;
        RECT 29.955 48.055 30.185 53.470 ;
        RECT 31.535 48.055 31.765 53.470 ;
        RECT 33.115 48.055 33.345 53.470 ;
        RECT 34.880 53.460 35.610 57.810 ;
        RECT 36.470 53.460 37.200 57.810 ;
        RECT 38.040 53.470 38.770 57.820 ;
        RECT 39.620 53.470 40.350 57.820 ;
        RECT 41.210 53.470 41.940 57.820 ;
        RECT 42.780 53.470 43.510 57.820 ;
        RECT 44.955 57.810 45.185 58.055 ;
        RECT 46.535 57.810 46.765 58.055 ;
        RECT 48.115 57.820 48.345 58.055 ;
        RECT 49.695 57.820 49.925 58.055 ;
        RECT 51.275 57.820 51.505 58.055 ;
        RECT 52.855 57.820 53.085 58.055 ;
        RECT 54.755 57.840 54.985 58.055 ;
        RECT 56.335 57.840 56.565 58.055 ;
        RECT 57.915 57.850 58.145 58.055 ;
        RECT 59.495 57.850 59.725 58.055 ;
        RECT 61.075 57.850 61.305 58.055 ;
        RECT 62.655 57.850 62.885 58.055 ;
        RECT 43.740 56.860 44.490 56.920 ;
        RECT 43.720 54.440 44.510 56.860 ;
        RECT 43.740 54.380 44.490 54.440 ;
        RECT 35.155 48.055 35.385 53.460 ;
        RECT 36.735 48.055 36.965 53.460 ;
        RECT 38.315 48.055 38.545 53.470 ;
        RECT 39.895 48.055 40.125 53.470 ;
        RECT 41.475 48.055 41.705 53.470 ;
        RECT 43.055 48.055 43.285 53.470 ;
        RECT 44.690 53.460 45.420 57.810 ;
        RECT 46.280 53.460 47.010 57.810 ;
        RECT 47.850 53.470 48.580 57.820 ;
        RECT 49.430 53.470 50.160 57.820 ;
        RECT 51.020 53.470 51.750 57.820 ;
        RECT 52.590 53.470 53.320 57.820 ;
        RECT 54.500 53.490 55.230 57.840 ;
        RECT 56.090 53.490 56.820 57.840 ;
        RECT 57.660 53.500 58.390 57.850 ;
        RECT 59.240 53.500 59.970 57.850 ;
        RECT 60.830 53.500 61.560 57.850 ;
        RECT 62.400 53.500 63.130 57.850 ;
        RECT 64.555 57.840 64.785 58.055 ;
        RECT 66.135 57.840 66.365 58.055 ;
        RECT 67.715 57.850 67.945 58.055 ;
        RECT 69.295 57.850 69.525 58.055 ;
        RECT 70.875 57.850 71.105 58.055 ;
        RECT 72.455 57.850 72.685 58.055 ;
        RECT 63.320 56.860 64.070 56.920 ;
        RECT 63.300 54.440 64.090 56.860 ;
        RECT 63.320 54.380 64.070 54.440 ;
        RECT 44.955 48.055 45.185 53.460 ;
        RECT 46.535 48.055 46.765 53.460 ;
        RECT 48.115 48.055 48.345 53.470 ;
        RECT 49.695 48.055 49.925 53.470 ;
        RECT 51.275 48.055 51.505 53.470 ;
        RECT 52.855 48.055 53.085 53.470 ;
        RECT 54.755 48.055 54.985 53.490 ;
        RECT 56.335 48.055 56.565 53.490 ;
        RECT 57.915 48.055 58.145 53.500 ;
        RECT 59.495 48.055 59.725 53.500 ;
        RECT 61.075 48.055 61.305 53.500 ;
        RECT 62.655 48.055 62.885 53.500 ;
        RECT 64.290 53.490 65.020 57.840 ;
        RECT 65.880 53.490 66.610 57.840 ;
        RECT 67.450 53.500 68.180 57.850 ;
        RECT 69.030 53.500 69.760 57.850 ;
        RECT 70.620 53.500 71.350 57.850 ;
        RECT 72.190 53.500 72.920 57.850 ;
        RECT 64.555 48.055 64.785 53.490 ;
        RECT 66.135 48.055 66.365 53.490 ;
        RECT 67.715 48.055 67.945 53.500 ;
        RECT 69.295 48.055 69.525 53.500 ;
        RECT 70.875 48.055 71.105 53.500 ;
        RECT 72.455 48.055 72.685 53.500 ;
        RECT 16.580 45.210 16.810 45.560 ;
        RECT 16.440 44.540 16.890 45.210 ;
        RECT 19.275 45.200 19.505 45.560 ;
        RECT 19.190 44.550 19.590 45.200 ;
        RECT 20.855 45.190 21.085 45.560 ;
        RECT 22.435 45.220 22.665 45.560 ;
        RECT 16.580 41.560 16.810 44.540 ;
        RECT 19.275 40.560 19.505 44.550 ;
        RECT 20.790 44.540 21.190 45.190 ;
        RECT 22.340 44.570 22.740 45.220 ;
        RECT 20.855 40.560 21.085 44.540 ;
        RECT 22.435 40.560 22.665 44.570 ;
        RECT 17.370 38.460 17.600 39.070 ;
        RECT 17.370 38.090 19.480 38.460 ;
        RECT 17.370 38.070 17.600 38.090 ;
        RECT 18.820 37.560 19.480 38.090 ;
        RECT 21.940 37.440 22.720 38.800 ;
        RECT 1.550 1.050 11.510 1.280 ;
      LAYER via ;
        RECT 22.135 103.175 22.505 103.545 ;
        RECT 16.490 96.620 16.840 97.290 ;
        RECT 19.240 96.630 19.540 97.280 ;
        RECT 20.840 96.640 21.140 97.290 ;
        RECT 22.390 96.610 22.690 97.260 ;
        RECT 1.620 84.640 11.610 85.240 ;
        RECT 14.980 84.340 15.280 84.990 ;
        RECT 16.560 84.330 16.860 84.980 ;
        RECT 18.150 84.330 18.450 84.980 ;
        RECT 19.730 84.330 20.030 84.980 ;
        RECT 21.310 84.330 21.610 84.980 ;
        RECT 22.900 84.330 23.200 84.980 ;
        RECT 25.000 84.020 25.630 88.370 ;
        RECT 26.590 84.020 27.220 88.370 ;
        RECT 28.160 84.010 28.790 88.360 ;
        RECT 29.740 84.010 30.370 88.360 ;
        RECT 31.330 84.010 31.960 88.360 ;
        RECT 32.900 84.010 33.530 88.360 ;
        RECT 34.930 84.020 35.560 88.370 ;
        RECT 36.520 84.020 37.150 88.370 ;
        RECT 38.090 84.010 38.720 88.360 ;
        RECT 39.670 84.010 40.300 88.360 ;
        RECT 41.260 84.010 41.890 88.360 ;
        RECT 42.830 84.010 43.460 88.360 ;
        RECT 43.770 84.970 44.460 87.390 ;
        RECT 44.740 84.020 45.370 88.370 ;
        RECT 46.330 84.020 46.960 88.370 ;
        RECT 47.900 84.010 48.530 88.360 ;
        RECT 49.480 84.010 50.110 88.360 ;
        RECT 51.070 84.010 51.700 88.360 ;
        RECT 52.640 84.010 53.270 88.360 ;
        RECT 54.550 83.990 55.180 88.340 ;
        RECT 56.140 83.990 56.770 88.340 ;
        RECT 57.710 83.980 58.340 88.330 ;
        RECT 59.290 83.980 59.920 88.330 ;
        RECT 60.880 83.980 61.510 88.330 ;
        RECT 62.450 83.980 63.080 88.330 ;
        RECT 63.350 84.970 64.040 87.390 ;
        RECT 64.340 83.990 64.970 88.340 ;
        RECT 65.930 83.990 66.560 88.340 ;
        RECT 67.500 83.980 68.130 88.330 ;
        RECT 69.080 83.980 69.710 88.330 ;
        RECT 70.670 83.980 71.300 88.330 ;
        RECT 72.240 83.980 72.870 88.330 ;
        RECT 25.010 72.970 25.640 77.320 ;
        RECT 26.600 72.970 27.230 77.320 ;
        RECT 28.170 72.960 28.800 77.310 ;
        RECT 29.750 72.960 30.380 77.310 ;
        RECT 31.340 72.960 31.970 77.310 ;
        RECT 32.910 72.960 33.540 77.310 ;
        RECT 33.900 73.840 34.590 76.260 ;
        RECT 34.940 72.970 35.570 77.320 ;
        RECT 36.530 72.970 37.160 77.320 ;
        RECT 38.100 72.960 38.730 77.310 ;
        RECT 39.680 72.960 40.310 77.310 ;
        RECT 41.270 72.960 41.900 77.310 ;
        RECT 42.840 72.960 43.470 77.310 ;
        RECT 44.750 72.970 45.380 77.320 ;
        RECT 46.340 72.970 46.970 77.320 ;
        RECT 47.910 72.960 48.540 77.310 ;
        RECT 49.490 72.960 50.120 77.310 ;
        RECT 51.080 72.960 51.710 77.310 ;
        RECT 52.650 72.960 53.280 77.310 ;
        RECT 53.570 73.850 54.260 76.270 ;
        RECT 54.560 72.940 55.190 77.290 ;
        RECT 56.150 72.940 56.780 77.290 ;
        RECT 57.720 72.930 58.350 77.280 ;
        RECT 59.300 72.930 59.930 77.280 ;
        RECT 60.890 72.930 61.520 77.280 ;
        RECT 62.460 72.930 63.090 77.280 ;
        RECT 64.350 72.940 64.980 77.290 ;
        RECT 65.940 72.940 66.570 77.290 ;
        RECT 67.510 72.930 68.140 77.280 ;
        RECT 69.090 72.930 69.720 77.280 ;
        RECT 70.680 72.930 71.310 77.280 ;
        RECT 72.250 72.930 72.880 77.280 ;
        RECT 25.010 64.510 25.640 68.860 ;
        RECT 26.600 64.510 27.230 68.860 ;
        RECT 28.170 64.520 28.800 68.870 ;
        RECT 29.750 64.520 30.380 68.870 ;
        RECT 31.340 64.520 31.970 68.870 ;
        RECT 32.910 64.520 33.540 68.870 ;
        RECT 33.900 65.570 34.590 67.990 ;
        RECT 17.695 62.030 17.955 62.880 ;
        RECT 19.275 62.030 19.535 62.880 ;
        RECT 19.935 62.030 20.355 62.880 ;
        RECT 20.775 62.030 21.035 62.880 ;
        RECT 22.345 62.030 22.605 62.880 ;
        RECT 2.565 60.805 2.825 61.425 ;
        RECT 3.525 60.805 3.785 61.425 ;
        RECT 4.485 60.805 4.745 61.425 ;
        RECT 5.445 60.805 5.705 61.425 ;
        RECT 6.405 60.805 6.665 61.425 ;
        RECT 7.365 60.805 7.625 61.425 ;
        RECT 7.925 60.805 8.205 61.425 ;
        RECT 8.505 60.805 8.765 61.425 ;
        RECT 9.465 60.805 9.725 61.425 ;
        RECT 10.425 60.805 10.685 61.425 ;
        RECT 11.385 60.805 11.645 61.425 ;
        RECT 12.345 60.805 12.605 61.425 ;
        RECT 13.305 60.805 13.565 61.425 ;
        RECT 34.940 64.510 35.570 68.860 ;
        RECT 36.530 64.510 37.160 68.860 ;
        RECT 38.100 64.520 38.730 68.870 ;
        RECT 39.680 64.520 40.310 68.870 ;
        RECT 41.270 64.520 41.900 68.870 ;
        RECT 42.840 64.520 43.470 68.870 ;
        RECT 44.750 64.510 45.380 68.860 ;
        RECT 46.340 64.510 46.970 68.860 ;
        RECT 47.910 64.520 48.540 68.870 ;
        RECT 49.490 64.520 50.120 68.870 ;
        RECT 51.080 64.520 51.710 68.870 ;
        RECT 52.650 64.520 53.280 68.870 ;
        RECT 53.570 65.560 54.260 67.980 ;
        RECT 54.560 64.540 55.190 68.890 ;
        RECT 56.150 64.540 56.780 68.890 ;
        RECT 57.720 64.550 58.350 68.900 ;
        RECT 59.300 64.550 59.930 68.900 ;
        RECT 60.890 64.550 61.520 68.900 ;
        RECT 62.460 64.550 63.090 68.900 ;
        RECT 64.350 64.540 64.980 68.890 ;
        RECT 65.940 64.540 66.570 68.890 ;
        RECT 67.510 64.550 68.140 68.900 ;
        RECT 69.090 64.550 69.720 68.900 ;
        RECT 70.680 64.550 71.310 68.900 ;
        RECT 72.250 64.550 72.880 68.900 ;
        RECT 1.530 56.730 11.530 57.200 ;
        RECT 14.980 56.840 15.280 57.490 ;
        RECT 16.560 56.850 16.860 57.500 ;
        RECT 18.150 56.850 18.450 57.500 ;
        RECT 19.730 56.850 20.030 57.500 ;
        RECT 21.310 56.850 21.610 57.500 ;
        RECT 22.900 56.850 23.200 57.500 ;
        RECT 25.000 53.460 25.630 57.810 ;
        RECT 26.590 53.460 27.220 57.810 ;
        RECT 28.160 53.470 28.790 57.820 ;
        RECT 29.740 53.470 30.370 57.820 ;
        RECT 31.330 53.470 31.960 57.820 ;
        RECT 32.900 53.470 33.530 57.820 ;
        RECT 34.930 53.460 35.560 57.810 ;
        RECT 36.520 53.460 37.150 57.810 ;
        RECT 38.090 53.470 38.720 57.820 ;
        RECT 39.670 53.470 40.300 57.820 ;
        RECT 41.260 53.470 41.890 57.820 ;
        RECT 42.830 53.470 43.460 57.820 ;
        RECT 43.770 54.440 44.460 56.860 ;
        RECT 44.740 53.460 45.370 57.810 ;
        RECT 46.330 53.460 46.960 57.810 ;
        RECT 47.900 53.470 48.530 57.820 ;
        RECT 49.480 53.470 50.110 57.820 ;
        RECT 51.070 53.470 51.700 57.820 ;
        RECT 52.640 53.470 53.270 57.820 ;
        RECT 54.550 53.490 55.180 57.840 ;
        RECT 56.140 53.490 56.770 57.840 ;
        RECT 57.710 53.500 58.340 57.850 ;
        RECT 59.290 53.500 59.920 57.850 ;
        RECT 60.880 53.500 61.510 57.850 ;
        RECT 62.450 53.500 63.080 57.850 ;
        RECT 63.350 54.440 64.040 56.860 ;
        RECT 64.340 53.490 64.970 57.840 ;
        RECT 65.930 53.490 66.560 57.840 ;
        RECT 67.500 53.500 68.130 57.850 ;
        RECT 69.080 53.500 69.710 57.850 ;
        RECT 70.670 53.500 71.300 57.850 ;
        RECT 72.240 53.500 72.870 57.850 ;
        RECT 16.490 44.540 16.840 45.210 ;
        RECT 19.240 44.550 19.540 45.200 ;
        RECT 20.840 44.540 21.140 45.190 ;
        RECT 22.390 44.570 22.690 45.220 ;
        RECT 22.135 38.285 22.505 38.655 ;
      LAYER met2 ;
        RECT 22.105 103.175 23.355 103.545 ;
        RECT 16.490 97.160 16.840 97.340 ;
        RECT 19.240 97.160 19.540 97.330 ;
        RECT 20.840 97.160 21.140 97.340 ;
        RECT 22.390 97.160 22.690 97.310 ;
        RECT 14.865 97.135 22.690 97.160 ;
        RECT 22.985 97.135 23.355 103.175 ;
        RECT 14.865 96.765 23.355 97.135 ;
        RECT 14.865 96.730 22.690 96.765 ;
        RECT 14.865 87.340 15.295 96.730 ;
        RECT 16.490 96.570 16.840 96.730 ;
        RECT 19.240 96.580 19.540 96.730 ;
        RECT 20.840 96.590 21.140 96.730 ;
        RECT 22.390 96.560 22.690 96.730 ;
        RECT 25.000 87.380 25.630 88.420 ;
        RECT 26.590 87.380 27.220 88.420 ;
        RECT 28.160 87.380 28.790 88.410 ;
        RECT 29.740 87.380 30.370 88.410 ;
        RECT 31.330 87.380 31.960 88.410 ;
        RECT 32.900 87.380 33.530 88.410 ;
        RECT 34.930 87.380 35.560 88.420 ;
        RECT 36.520 87.380 37.150 88.420 ;
        RECT 38.090 87.380 38.720 88.410 ;
        RECT 39.670 87.380 40.300 88.410 ;
        RECT 41.260 87.380 41.890 88.410 ;
        RECT 42.830 87.380 43.460 88.410 ;
        RECT 43.770 87.380 44.460 87.440 ;
        RECT 44.740 87.380 45.370 88.420 ;
        RECT 46.330 87.380 46.960 88.420 ;
        RECT 47.900 87.380 48.530 88.410 ;
        RECT 49.480 87.380 50.110 88.410 ;
        RECT 51.070 87.380 51.700 88.410 ;
        RECT 52.640 87.380 53.270 88.410 ;
        RECT 54.550 87.380 55.180 88.390 ;
        RECT 56.140 87.380 56.770 88.390 ;
        RECT 57.710 87.380 58.340 88.380 ;
        RECT 59.290 87.380 59.920 88.380 ;
        RECT 60.880 87.380 61.510 88.380 ;
        RECT 62.450 87.380 63.080 88.380 ;
        RECT 63.350 87.380 64.040 87.440 ;
        RECT 64.340 87.380 64.970 88.390 ;
        RECT 65.930 87.380 66.560 88.390 ;
        RECT 67.500 87.380 68.130 88.380 ;
        RECT 69.080 87.380 69.710 88.380 ;
        RECT 70.670 87.380 71.300 88.380 ;
        RECT 72.240 87.380 72.870 88.380 ;
        RECT 25.000 87.340 72.870 87.380 ;
        RECT 1.600 84.950 72.870 87.340 ;
        RECT 1.600 84.260 25.630 84.950 ;
        RECT 14.865 84.255 15.295 84.260 ;
        RECT 25.000 83.970 25.630 84.260 ;
        RECT 26.590 83.970 27.220 84.950 ;
        RECT 28.160 83.960 28.790 84.950 ;
        RECT 29.740 83.960 30.370 84.950 ;
        RECT 31.330 83.960 31.960 84.950 ;
        RECT 32.900 83.960 33.530 84.950 ;
        RECT 34.930 83.970 35.560 84.950 ;
        RECT 36.520 83.970 37.150 84.950 ;
        RECT 38.090 83.960 38.720 84.950 ;
        RECT 39.670 83.960 40.300 84.950 ;
        RECT 41.260 83.960 41.890 84.950 ;
        RECT 42.830 83.960 43.460 84.950 ;
        RECT 43.770 84.920 44.460 84.950 ;
        RECT 44.740 83.970 45.370 84.950 ;
        RECT 46.330 83.970 46.960 84.950 ;
        RECT 47.900 83.960 48.530 84.950 ;
        RECT 49.480 83.960 50.110 84.950 ;
        RECT 51.070 83.960 51.700 84.950 ;
        RECT 52.640 83.960 53.270 84.950 ;
        RECT 54.550 83.940 55.180 84.950 ;
        RECT 56.140 83.940 56.770 84.950 ;
        RECT 57.710 83.930 58.340 84.950 ;
        RECT 59.290 83.930 59.920 84.950 ;
        RECT 60.880 83.930 61.510 84.950 ;
        RECT 62.450 83.930 63.080 84.950 ;
        RECT 63.350 84.920 64.040 84.950 ;
        RECT 64.340 83.940 64.970 84.950 ;
        RECT 65.930 83.940 66.560 84.950 ;
        RECT 67.500 83.930 68.130 84.950 ;
        RECT 69.080 83.930 69.710 84.950 ;
        RECT 70.670 83.930 71.300 84.950 ;
        RECT 72.240 83.930 72.870 84.950 ;
        RECT 25.010 76.270 25.640 77.370 ;
        RECT 26.600 76.270 27.230 77.370 ;
        RECT 28.170 76.270 28.800 77.360 ;
        RECT 29.750 76.270 30.380 77.360 ;
        RECT 31.340 76.270 31.970 77.360 ;
        RECT 32.910 76.270 33.540 77.360 ;
        RECT 33.900 76.270 34.590 76.310 ;
        RECT 34.940 76.270 35.570 77.370 ;
        RECT 36.530 76.270 37.160 77.370 ;
        RECT 38.100 76.270 38.730 77.360 ;
        RECT 39.680 76.270 40.310 77.360 ;
        RECT 41.270 76.270 41.900 77.360 ;
        RECT 42.840 76.270 43.470 77.360 ;
        RECT 44.750 76.270 45.380 77.370 ;
        RECT 46.340 76.270 46.970 77.370 ;
        RECT 47.910 76.270 48.540 77.360 ;
        RECT 49.490 76.270 50.120 77.360 ;
        RECT 51.080 76.270 51.710 77.360 ;
        RECT 52.650 76.270 53.280 77.360 ;
        RECT 53.570 76.270 54.260 76.320 ;
        RECT 54.560 76.270 55.190 77.340 ;
        RECT 56.150 76.270 56.780 77.340 ;
        RECT 57.720 76.270 58.350 77.330 ;
        RECT 59.300 76.270 59.930 77.330 ;
        RECT 60.890 76.270 61.520 77.330 ;
        RECT 62.460 76.270 63.090 77.330 ;
        RECT 64.350 76.270 64.980 77.340 ;
        RECT 65.940 76.270 66.570 77.340 ;
        RECT 67.510 76.270 68.140 77.330 ;
        RECT 69.090 76.270 69.720 77.330 ;
        RECT 70.680 76.270 71.310 77.330 ;
        RECT 72.250 76.270 72.880 77.330 ;
        RECT 25.010 73.840 72.880 76.270 ;
        RECT 25.010 72.920 25.640 73.840 ;
        RECT 26.600 72.920 27.230 73.840 ;
        RECT 28.170 72.910 28.800 73.840 ;
        RECT 29.750 72.910 30.380 73.840 ;
        RECT 31.340 72.910 31.970 73.840 ;
        RECT 32.910 72.910 33.540 73.840 ;
        RECT 33.900 73.790 34.590 73.840 ;
        RECT 34.940 72.920 35.570 73.840 ;
        RECT 36.530 72.920 37.160 73.840 ;
        RECT 38.100 72.910 38.730 73.840 ;
        RECT 39.680 72.910 40.310 73.840 ;
        RECT 41.270 72.910 41.900 73.840 ;
        RECT 42.840 72.910 43.470 73.840 ;
        RECT 44.750 72.920 45.380 73.840 ;
        RECT 46.340 72.920 46.970 73.840 ;
        RECT 47.910 72.910 48.540 73.840 ;
        RECT 49.490 72.910 50.120 73.840 ;
        RECT 51.080 72.910 51.710 73.840 ;
        RECT 52.650 72.910 53.280 73.840 ;
        RECT 53.570 73.800 54.260 73.840 ;
        RECT 54.560 72.890 55.190 73.840 ;
        RECT 56.150 72.890 56.780 73.840 ;
        RECT 57.720 72.880 58.350 73.840 ;
        RECT 59.300 72.880 59.930 73.840 ;
        RECT 60.890 72.880 61.520 73.840 ;
        RECT 62.460 72.880 63.090 73.840 ;
        RECT 64.350 72.890 64.980 73.840 ;
        RECT 65.940 72.890 66.570 73.840 ;
        RECT 67.510 72.880 68.140 73.840 ;
        RECT 69.090 72.880 69.720 73.840 ;
        RECT 70.680 72.880 71.310 73.840 ;
        RECT 72.250 72.880 72.880 73.840 ;
        RECT 25.010 67.990 25.640 68.910 ;
        RECT 26.600 67.990 27.230 68.910 ;
        RECT 28.170 67.990 28.800 68.920 ;
        RECT 29.750 67.990 30.380 68.920 ;
        RECT 31.340 67.990 31.970 68.920 ;
        RECT 32.910 67.990 33.540 68.920 ;
        RECT 33.900 67.990 34.590 68.040 ;
        RECT 34.940 67.990 35.570 68.910 ;
        RECT 36.530 67.990 37.160 68.910 ;
        RECT 38.100 67.990 38.730 68.920 ;
        RECT 39.680 67.990 40.310 68.920 ;
        RECT 41.270 67.990 41.900 68.920 ;
        RECT 42.840 67.990 43.470 68.920 ;
        RECT 44.750 67.990 45.380 68.910 ;
        RECT 46.340 67.990 46.970 68.910 ;
        RECT 47.910 67.990 48.540 68.920 ;
        RECT 49.490 67.990 50.120 68.920 ;
        RECT 51.080 67.990 51.710 68.920 ;
        RECT 52.650 67.990 53.280 68.920 ;
        RECT 53.570 67.990 54.260 68.030 ;
        RECT 54.560 67.990 55.190 68.940 ;
        RECT 56.150 67.990 56.780 68.940 ;
        RECT 57.720 67.990 58.350 68.950 ;
        RECT 59.300 67.990 59.930 68.950 ;
        RECT 60.890 67.990 61.520 68.950 ;
        RECT 62.460 67.990 63.090 68.950 ;
        RECT 64.350 67.990 64.980 68.940 ;
        RECT 65.940 67.990 66.570 68.940 ;
        RECT 67.510 67.990 68.140 68.950 ;
        RECT 69.090 67.990 69.720 68.950 ;
        RECT 70.680 67.990 71.310 68.950 ;
        RECT 72.250 67.990 72.880 68.950 ;
        RECT 25.010 65.560 72.880 67.990 ;
        RECT 25.010 64.460 25.640 65.560 ;
        RECT 26.600 64.460 27.230 65.560 ;
        RECT 28.170 64.470 28.800 65.560 ;
        RECT 29.750 64.470 30.380 65.560 ;
        RECT 31.340 64.470 31.970 65.560 ;
        RECT 32.910 64.470 33.540 65.560 ;
        RECT 33.900 65.520 34.590 65.560 ;
        RECT 34.940 64.460 35.570 65.560 ;
        RECT 36.530 64.460 37.160 65.560 ;
        RECT 38.100 64.470 38.730 65.560 ;
        RECT 39.680 64.470 40.310 65.560 ;
        RECT 41.270 64.470 41.900 65.560 ;
        RECT 42.840 64.470 43.470 65.560 ;
        RECT 44.750 64.460 45.380 65.560 ;
        RECT 46.340 64.460 46.970 65.560 ;
        RECT 47.910 64.470 48.540 65.560 ;
        RECT 49.490 64.470 50.120 65.560 ;
        RECT 51.080 64.470 51.710 65.560 ;
        RECT 52.650 64.470 53.280 65.560 ;
        RECT 53.570 65.510 54.260 65.560 ;
        RECT 54.560 64.490 55.190 65.560 ;
        RECT 56.150 64.490 56.780 65.560 ;
        RECT 57.720 64.500 58.350 65.560 ;
        RECT 59.300 64.500 59.930 65.560 ;
        RECT 60.890 64.500 61.520 65.560 ;
        RECT 62.460 64.500 63.090 65.560 ;
        RECT 64.350 64.490 64.980 65.560 ;
        RECT 65.940 64.490 66.570 65.560 ;
        RECT 67.510 64.500 68.140 65.560 ;
        RECT 69.090 64.500 69.720 65.560 ;
        RECT 70.680 64.500 71.310 65.560 ;
        RECT 72.250 64.500 72.880 65.560 ;
        RECT 17.695 62.880 17.955 62.930 ;
        RECT 19.275 62.880 19.535 62.930 ;
        RECT 19.935 62.880 20.355 62.930 ;
        RECT 20.775 62.880 21.035 62.930 ;
        RECT 22.345 62.880 22.605 62.930 ;
        RECT 17.695 62.680 22.605 62.880 ;
        RECT 15.580 62.060 25.040 62.680 ;
        RECT 2.565 61.425 2.825 61.475 ;
        RECT 3.525 61.425 3.785 61.475 ;
        RECT 4.485 61.425 4.745 61.475 ;
        RECT 5.445 61.425 5.705 61.475 ;
        RECT 6.405 61.425 6.665 61.475 ;
        RECT 7.365 61.425 7.625 61.485 ;
        RECT 7.925 61.425 8.205 61.475 ;
        RECT 8.505 61.425 8.765 61.475 ;
        RECT 9.465 61.425 9.725 61.475 ;
        RECT 10.425 61.425 10.685 61.475 ;
        RECT 11.385 61.425 11.645 61.475 ;
        RECT 12.345 61.425 12.605 61.475 ;
        RECT 13.305 61.430 13.565 61.475 ;
        RECT 15.580 61.430 16.200 62.060 ;
        RECT 17.695 62.030 22.605 62.060 ;
        RECT 17.695 61.980 17.955 62.030 ;
        RECT 19.275 61.980 19.535 62.030 ;
        RECT 19.935 61.980 20.355 62.030 ;
        RECT 20.775 61.980 21.035 62.030 ;
        RECT 22.345 61.980 22.605 62.030 ;
        RECT 13.305 61.425 16.200 61.430 ;
        RECT 2.565 60.810 16.200 61.425 ;
        RECT 2.565 60.805 13.565 60.810 ;
        RECT 2.565 60.755 2.825 60.805 ;
        RECT 3.525 60.755 3.785 60.805 ;
        RECT 4.485 60.755 4.745 60.805 ;
        RECT 5.445 60.755 5.705 60.805 ;
        RECT 6.405 60.755 6.665 60.805 ;
        RECT 7.365 60.765 7.625 60.805 ;
        RECT 7.925 60.755 8.205 60.805 ;
        RECT 8.505 60.755 8.765 60.805 ;
        RECT 9.465 60.755 9.725 60.805 ;
        RECT 10.425 60.755 10.685 60.805 ;
        RECT 11.385 60.755 11.645 60.805 ;
        RECT 12.345 60.755 12.605 60.805 ;
        RECT 13.305 60.755 13.565 60.805 ;
        RECT 24.420 57.860 25.040 62.060 ;
        RECT 24.420 57.700 25.630 57.860 ;
        RECT 1.490 56.880 25.630 57.700 ;
        RECT 26.590 56.880 27.220 57.860 ;
        RECT 28.160 56.880 28.790 57.870 ;
        RECT 29.740 56.880 30.370 57.870 ;
        RECT 31.330 56.880 31.960 57.870 ;
        RECT 32.900 56.880 33.530 57.870 ;
        RECT 34.930 56.880 35.560 57.860 ;
        RECT 36.520 56.880 37.150 57.860 ;
        RECT 38.090 56.880 38.720 57.870 ;
        RECT 39.670 56.880 40.300 57.870 ;
        RECT 41.260 56.880 41.890 57.870 ;
        RECT 42.830 56.880 43.460 57.870 ;
        RECT 43.770 56.880 44.460 56.910 ;
        RECT 44.740 56.880 45.370 57.860 ;
        RECT 46.330 56.880 46.960 57.860 ;
        RECT 47.900 56.880 48.530 57.870 ;
        RECT 49.480 56.880 50.110 57.870 ;
        RECT 51.070 56.880 51.700 57.870 ;
        RECT 52.640 56.880 53.270 57.870 ;
        RECT 54.550 56.880 55.180 57.890 ;
        RECT 56.140 56.880 56.770 57.890 ;
        RECT 57.710 56.880 58.340 57.900 ;
        RECT 59.290 56.880 59.920 57.900 ;
        RECT 60.880 56.880 61.510 57.900 ;
        RECT 62.450 56.880 63.080 57.900 ;
        RECT 63.350 56.880 64.040 56.910 ;
        RECT 64.340 56.880 64.970 57.890 ;
        RECT 65.930 56.880 66.560 57.890 ;
        RECT 67.500 56.880 68.130 57.900 ;
        RECT 69.080 56.880 69.710 57.900 ;
        RECT 70.670 56.880 71.300 57.900 ;
        RECT 72.240 56.880 72.870 57.900 ;
        RECT 1.490 55.760 72.870 56.880 ;
        RECT 14.865 45.100 15.295 55.760 ;
        RECT 25.000 54.450 72.870 55.760 ;
        RECT 25.000 53.410 25.630 54.450 ;
        RECT 26.590 53.410 27.220 54.450 ;
        RECT 28.160 53.420 28.790 54.450 ;
        RECT 29.740 53.420 30.370 54.450 ;
        RECT 31.330 53.420 31.960 54.450 ;
        RECT 32.900 53.420 33.530 54.450 ;
        RECT 34.930 53.410 35.560 54.450 ;
        RECT 36.520 53.410 37.150 54.450 ;
        RECT 38.090 53.420 38.720 54.450 ;
        RECT 39.670 53.420 40.300 54.450 ;
        RECT 41.260 53.420 41.890 54.450 ;
        RECT 42.830 53.420 43.460 54.450 ;
        RECT 43.770 54.390 44.460 54.450 ;
        RECT 44.740 53.410 45.370 54.450 ;
        RECT 46.330 53.410 46.960 54.450 ;
        RECT 47.900 53.420 48.530 54.450 ;
        RECT 49.480 53.420 50.110 54.450 ;
        RECT 51.070 53.420 51.700 54.450 ;
        RECT 52.640 53.420 53.270 54.450 ;
        RECT 54.550 53.440 55.180 54.450 ;
        RECT 56.140 53.440 56.770 54.450 ;
        RECT 57.710 53.450 58.340 54.450 ;
        RECT 59.290 53.450 59.920 54.450 ;
        RECT 60.880 53.450 61.510 54.450 ;
        RECT 62.450 53.450 63.080 54.450 ;
        RECT 63.350 54.390 64.040 54.450 ;
        RECT 64.340 53.440 64.970 54.450 ;
        RECT 65.930 53.440 66.560 54.450 ;
        RECT 67.500 53.450 68.130 54.450 ;
        RECT 69.080 53.450 69.710 54.450 ;
        RECT 70.670 53.450 71.300 54.450 ;
        RECT 72.240 53.450 72.870 54.450 ;
        RECT 16.490 45.100 16.840 45.260 ;
        RECT 19.240 45.100 19.540 45.250 ;
        RECT 20.840 45.100 21.140 45.240 ;
        RECT 22.390 45.100 22.690 45.270 ;
        RECT 14.865 45.065 22.690 45.100 ;
        RECT 14.865 44.695 23.355 45.065 ;
        RECT 14.865 44.670 22.690 44.695 ;
        RECT 16.490 44.490 16.840 44.670 ;
        RECT 19.240 44.500 19.540 44.670 ;
        RECT 20.840 44.490 21.140 44.670 ;
        RECT 22.390 44.520 22.690 44.670 ;
        RECT 22.985 38.655 23.355 44.695 ;
        RECT 22.105 38.285 23.355 38.655 ;
      LAYER via2 ;
        RECT 43.660 85.040 59.820 86.610 ;
        RECT 43.750 74.300 59.880 75.870 ;
        RECT 43.750 65.960 59.880 67.530 ;
        RECT 43.660 55.220 59.820 56.790 ;
      LAYER met3 ;
        RECT 43.600 109.230 60.220 133.480 ;
        RECT 43.600 105.230 60.260 109.230 ;
        RECT 43.640 86.660 60.260 105.230 ;
        RECT 43.620 74.160 60.260 86.660 ;
        RECT 43.620 67.670 60.240 74.160 ;
        RECT 43.620 60.100 60.260 67.670 ;
        RECT 43.620 55.170 60.310 60.100 ;
        RECT 43.690 8.600 60.310 55.170 ;
      LAYER via3 ;
        RECT 44.270 9.340 59.430 66.680 ;
      LAYER met4 ;
        RECT 0.460 46.870 72.360 67.320 ;
        RECT 0.270 41.070 72.360 46.870 ;
        RECT 0.460 1.300 72.360 41.070 ;
      LAYER via4 ;
        RECT 0.270 41.070 72.240 46.870 ;
      LAYER met5 ;
        RECT 0.150 40.950 72.360 46.990 ;
    END
  END vss
  OBS
      LAYER li1 ;
        RECT 15.285 140.585 15.785 140.755 ;
        RECT 16.075 140.585 16.575 140.755 ;
        RECT 16.865 140.585 17.365 140.755 ;
        RECT 17.655 140.585 18.155 140.755 ;
        RECT 18.445 140.585 18.945 140.755 ;
        RECT 19.235 140.585 19.735 140.755 ;
        RECT 20.025 140.585 20.525 140.755 ;
        RECT 20.815 140.585 21.315 140.755 ;
        RECT 21.605 140.585 22.105 140.755 ;
        RECT 22.395 140.585 22.895 140.755 ;
        RECT 25.470 140.580 25.970 140.750 ;
        RECT 26.260 140.580 26.760 140.750 ;
        RECT 27.050 140.580 27.550 140.750 ;
        RECT 27.840 140.580 28.340 140.750 ;
        RECT 28.630 140.580 29.130 140.750 ;
        RECT 29.420 140.580 29.920 140.750 ;
        RECT 30.210 140.580 30.710 140.750 ;
        RECT 31.000 140.580 31.500 140.750 ;
        RECT 31.790 140.580 32.290 140.750 ;
        RECT 32.580 140.580 33.080 140.750 ;
        RECT 35.410 140.580 35.910 140.750 ;
        RECT 36.200 140.580 36.700 140.750 ;
        RECT 36.990 140.580 37.490 140.750 ;
        RECT 37.780 140.580 38.280 140.750 ;
        RECT 38.570 140.580 39.070 140.750 ;
        RECT 39.360 140.580 39.860 140.750 ;
        RECT 40.150 140.580 40.650 140.750 ;
        RECT 40.940 140.580 41.440 140.750 ;
        RECT 41.730 140.580 42.230 140.750 ;
        RECT 42.520 140.580 43.020 140.750 ;
        RECT 45.210 140.580 45.710 140.750 ;
        RECT 46.000 140.580 46.500 140.750 ;
        RECT 46.790 140.580 47.290 140.750 ;
        RECT 47.580 140.580 48.080 140.750 ;
        RECT 48.370 140.580 48.870 140.750 ;
        RECT 49.160 140.580 49.660 140.750 ;
        RECT 49.950 140.580 50.450 140.750 ;
        RECT 50.740 140.580 51.240 140.750 ;
        RECT 51.530 140.580 52.030 140.750 ;
        RECT 52.320 140.580 52.820 140.750 ;
        RECT 55.010 140.580 55.510 140.750 ;
        RECT 55.800 140.580 56.300 140.750 ;
        RECT 56.590 140.580 57.090 140.750 ;
        RECT 57.380 140.580 57.880 140.750 ;
        RECT 58.170 140.580 58.670 140.750 ;
        RECT 58.960 140.580 59.460 140.750 ;
        RECT 59.750 140.580 60.250 140.750 ;
        RECT 60.540 140.580 61.040 140.750 ;
        RECT 61.330 140.580 61.830 140.750 ;
        RECT 62.120 140.580 62.620 140.750 ;
        RECT 64.810 140.580 65.310 140.750 ;
        RECT 65.600 140.580 66.100 140.750 ;
        RECT 66.390 140.580 66.890 140.750 ;
        RECT 67.180 140.580 67.680 140.750 ;
        RECT 67.970 140.580 68.470 140.750 ;
        RECT 68.760 140.580 69.260 140.750 ;
        RECT 69.550 140.580 70.050 140.750 ;
        RECT 70.340 140.580 70.840 140.750 ;
        RECT 71.130 140.580 71.630 140.750 ;
        RECT 71.920 140.580 72.420 140.750 ;
        RECT 15.845 130.325 16.015 140.365 ;
        RECT 17.425 130.325 17.595 140.365 ;
        RECT 19.005 130.325 19.175 140.365 ;
        RECT 20.585 130.325 20.755 140.365 ;
        RECT 22.165 130.325 22.335 140.365 ;
        RECT 15.285 129.935 15.785 130.105 ;
        RECT 16.075 129.935 16.575 130.105 ;
        RECT 16.865 129.935 17.365 130.105 ;
        RECT 17.655 129.935 18.155 130.105 ;
        RECT 18.445 129.935 18.945 130.105 ;
        RECT 19.235 129.935 19.735 130.105 ;
        RECT 20.025 129.935 20.525 130.105 ;
        RECT 20.815 129.935 21.315 130.105 ;
        RECT 21.605 129.935 22.105 130.105 ;
        RECT 22.395 129.935 22.895 130.105 ;
        RECT 25.470 129.940 25.970 130.110 ;
        RECT 26.260 129.940 26.760 130.110 ;
        RECT 27.050 129.940 27.550 130.110 ;
        RECT 27.840 129.940 28.340 130.110 ;
        RECT 28.630 129.940 29.130 130.110 ;
        RECT 29.420 129.940 29.920 130.110 ;
        RECT 30.210 129.940 30.710 130.110 ;
        RECT 31.000 129.940 31.500 130.110 ;
        RECT 31.790 129.940 32.290 130.110 ;
        RECT 32.580 129.940 33.080 130.110 ;
        RECT 35.410 129.940 35.910 130.110 ;
        RECT 36.200 129.940 36.700 130.110 ;
        RECT 36.990 129.940 37.490 130.110 ;
        RECT 37.780 129.940 38.280 130.110 ;
        RECT 38.570 129.940 39.070 130.110 ;
        RECT 39.360 129.940 39.860 130.110 ;
        RECT 40.150 129.940 40.650 130.110 ;
        RECT 40.940 129.940 41.440 130.110 ;
        RECT 41.730 129.940 42.230 130.110 ;
        RECT 42.520 129.940 43.020 130.110 ;
        RECT 45.210 129.940 45.710 130.110 ;
        RECT 46.000 129.940 46.500 130.110 ;
        RECT 46.790 129.940 47.290 130.110 ;
        RECT 47.580 129.940 48.080 130.110 ;
        RECT 48.370 129.940 48.870 130.110 ;
        RECT 49.160 129.940 49.660 130.110 ;
        RECT 49.950 129.940 50.450 130.110 ;
        RECT 50.740 129.940 51.240 130.110 ;
        RECT 51.530 129.940 52.030 130.110 ;
        RECT 52.320 129.940 52.820 130.110 ;
        RECT 55.010 129.940 55.510 130.110 ;
        RECT 55.800 129.940 56.300 130.110 ;
        RECT 56.590 129.940 57.090 130.110 ;
        RECT 57.380 129.940 57.880 130.110 ;
        RECT 58.170 129.940 58.670 130.110 ;
        RECT 58.960 129.940 59.460 130.110 ;
        RECT 59.750 129.940 60.250 130.110 ;
        RECT 60.540 129.940 61.040 130.110 ;
        RECT 61.330 129.940 61.830 130.110 ;
        RECT 62.120 129.940 62.620 130.110 ;
        RECT 64.810 129.940 65.310 130.110 ;
        RECT 65.600 129.940 66.100 130.110 ;
        RECT 66.390 129.940 66.890 130.110 ;
        RECT 67.180 129.940 67.680 130.110 ;
        RECT 67.970 129.940 68.470 130.110 ;
        RECT 68.760 129.940 69.260 130.110 ;
        RECT 69.550 129.940 70.050 130.110 ;
        RECT 70.340 129.940 70.840 130.110 ;
        RECT 71.130 129.940 71.630 130.110 ;
        RECT 71.920 129.940 72.420 130.110 ;
        RECT 15.285 129.405 15.785 129.575 ;
        RECT 16.075 129.405 16.575 129.575 ;
        RECT 16.865 129.405 17.365 129.575 ;
        RECT 17.655 129.405 18.155 129.575 ;
        RECT 18.445 129.405 18.945 129.575 ;
        RECT 19.235 129.405 19.735 129.575 ;
        RECT 20.025 129.405 20.525 129.575 ;
        RECT 20.815 129.405 21.315 129.575 ;
        RECT 21.605 129.405 22.105 129.575 ;
        RECT 22.395 129.405 22.895 129.575 ;
        RECT 25.470 129.400 25.970 129.570 ;
        RECT 26.260 129.400 26.760 129.570 ;
        RECT 27.050 129.400 27.550 129.570 ;
        RECT 27.840 129.400 28.340 129.570 ;
        RECT 28.630 129.400 29.130 129.570 ;
        RECT 29.420 129.400 29.920 129.570 ;
        RECT 30.210 129.400 30.710 129.570 ;
        RECT 31.000 129.400 31.500 129.570 ;
        RECT 31.790 129.400 32.290 129.570 ;
        RECT 32.580 129.400 33.080 129.570 ;
        RECT 35.410 129.400 35.910 129.570 ;
        RECT 36.200 129.400 36.700 129.570 ;
        RECT 36.990 129.400 37.490 129.570 ;
        RECT 37.780 129.400 38.280 129.570 ;
        RECT 38.570 129.400 39.070 129.570 ;
        RECT 39.360 129.400 39.860 129.570 ;
        RECT 40.150 129.400 40.650 129.570 ;
        RECT 40.940 129.400 41.440 129.570 ;
        RECT 41.730 129.400 42.230 129.570 ;
        RECT 42.520 129.400 43.020 129.570 ;
        RECT 45.210 129.400 45.710 129.570 ;
        RECT 46.000 129.400 46.500 129.570 ;
        RECT 46.790 129.400 47.290 129.570 ;
        RECT 47.580 129.400 48.080 129.570 ;
        RECT 48.370 129.400 48.870 129.570 ;
        RECT 49.160 129.400 49.660 129.570 ;
        RECT 49.950 129.400 50.450 129.570 ;
        RECT 50.740 129.400 51.240 129.570 ;
        RECT 51.530 129.400 52.030 129.570 ;
        RECT 52.320 129.400 52.820 129.570 ;
        RECT 55.010 129.400 55.510 129.570 ;
        RECT 55.800 129.400 56.300 129.570 ;
        RECT 56.590 129.400 57.090 129.570 ;
        RECT 57.380 129.400 57.880 129.570 ;
        RECT 58.170 129.400 58.670 129.570 ;
        RECT 58.960 129.400 59.460 129.570 ;
        RECT 59.750 129.400 60.250 129.570 ;
        RECT 60.540 129.400 61.040 129.570 ;
        RECT 61.330 129.400 61.830 129.570 ;
        RECT 62.120 129.400 62.620 129.570 ;
        RECT 64.810 129.400 65.310 129.570 ;
        RECT 65.600 129.400 66.100 129.570 ;
        RECT 66.390 129.400 66.890 129.570 ;
        RECT 67.180 129.400 67.680 129.570 ;
        RECT 67.970 129.400 68.470 129.570 ;
        RECT 68.760 129.400 69.260 129.570 ;
        RECT 69.550 129.400 70.050 129.570 ;
        RECT 70.340 129.400 70.840 129.570 ;
        RECT 71.130 129.400 71.630 129.570 ;
        RECT 71.920 129.400 72.420 129.570 ;
        RECT 15.845 119.145 16.015 129.185 ;
        RECT 17.425 119.145 17.595 129.185 ;
        RECT 19.005 119.145 19.175 129.185 ;
        RECT 20.585 119.145 20.755 129.185 ;
        RECT 22.165 119.145 22.335 129.185 ;
        RECT 15.285 118.755 15.785 118.925 ;
        RECT 16.075 118.755 16.575 118.925 ;
        RECT 16.865 118.755 17.365 118.925 ;
        RECT 17.655 118.755 18.155 118.925 ;
        RECT 18.445 118.755 18.945 118.925 ;
        RECT 19.235 118.755 19.735 118.925 ;
        RECT 20.025 118.755 20.525 118.925 ;
        RECT 20.815 118.755 21.315 118.925 ;
        RECT 21.605 118.755 22.105 118.925 ;
        RECT 22.395 118.755 22.895 118.925 ;
        RECT 25.470 118.760 25.970 118.930 ;
        RECT 26.260 118.760 26.760 118.930 ;
        RECT 27.050 118.760 27.550 118.930 ;
        RECT 27.840 118.760 28.340 118.930 ;
        RECT 28.630 118.760 29.130 118.930 ;
        RECT 29.420 118.760 29.920 118.930 ;
        RECT 30.210 118.760 30.710 118.930 ;
        RECT 31.000 118.760 31.500 118.930 ;
        RECT 31.790 118.760 32.290 118.930 ;
        RECT 32.580 118.760 33.080 118.930 ;
        RECT 35.410 118.760 35.910 118.930 ;
        RECT 36.200 118.760 36.700 118.930 ;
        RECT 36.990 118.760 37.490 118.930 ;
        RECT 37.780 118.760 38.280 118.930 ;
        RECT 38.570 118.760 39.070 118.930 ;
        RECT 39.360 118.760 39.860 118.930 ;
        RECT 40.150 118.760 40.650 118.930 ;
        RECT 40.940 118.760 41.440 118.930 ;
        RECT 41.730 118.760 42.230 118.930 ;
        RECT 42.520 118.760 43.020 118.930 ;
        RECT 45.210 118.760 45.710 118.930 ;
        RECT 46.000 118.760 46.500 118.930 ;
        RECT 46.790 118.760 47.290 118.930 ;
        RECT 47.580 118.760 48.080 118.930 ;
        RECT 48.370 118.760 48.870 118.930 ;
        RECT 49.160 118.760 49.660 118.930 ;
        RECT 49.950 118.760 50.450 118.930 ;
        RECT 50.740 118.760 51.240 118.930 ;
        RECT 51.530 118.760 52.030 118.930 ;
        RECT 52.320 118.760 52.820 118.930 ;
        RECT 55.010 118.760 55.510 118.930 ;
        RECT 55.800 118.760 56.300 118.930 ;
        RECT 56.590 118.760 57.090 118.930 ;
        RECT 57.380 118.760 57.880 118.930 ;
        RECT 58.170 118.760 58.670 118.930 ;
        RECT 58.960 118.760 59.460 118.930 ;
        RECT 59.750 118.760 60.250 118.930 ;
        RECT 60.540 118.760 61.040 118.930 ;
        RECT 61.330 118.760 61.830 118.930 ;
        RECT 62.120 118.760 62.620 118.930 ;
        RECT 64.810 118.760 65.310 118.930 ;
        RECT 65.600 118.760 66.100 118.930 ;
        RECT 66.390 118.760 66.890 118.930 ;
        RECT 67.180 118.760 67.680 118.930 ;
        RECT 67.970 118.760 68.470 118.930 ;
        RECT 68.760 118.760 69.260 118.930 ;
        RECT 69.550 118.760 70.050 118.930 ;
        RECT 70.340 118.760 70.840 118.930 ;
        RECT 71.130 118.760 71.630 118.930 ;
        RECT 71.920 118.760 72.420 118.930 ;
        RECT 25.470 118.220 25.970 118.390 ;
        RECT 26.260 118.220 26.760 118.390 ;
        RECT 27.050 118.220 27.550 118.390 ;
        RECT 27.840 118.220 28.340 118.390 ;
        RECT 28.630 118.220 29.130 118.390 ;
        RECT 29.420 118.220 29.920 118.390 ;
        RECT 30.210 118.220 30.710 118.390 ;
        RECT 31.000 118.220 31.500 118.390 ;
        RECT 31.790 118.220 32.290 118.390 ;
        RECT 32.580 118.220 33.080 118.390 ;
        RECT 35.410 118.220 35.910 118.390 ;
        RECT 36.200 118.220 36.700 118.390 ;
        RECT 36.990 118.220 37.490 118.390 ;
        RECT 37.780 118.220 38.280 118.390 ;
        RECT 38.570 118.220 39.070 118.390 ;
        RECT 39.360 118.220 39.860 118.390 ;
        RECT 40.150 118.220 40.650 118.390 ;
        RECT 40.940 118.220 41.440 118.390 ;
        RECT 41.730 118.220 42.230 118.390 ;
        RECT 42.520 118.220 43.020 118.390 ;
        RECT 45.210 118.220 45.710 118.390 ;
        RECT 46.000 118.220 46.500 118.390 ;
        RECT 46.790 118.220 47.290 118.390 ;
        RECT 47.580 118.220 48.080 118.390 ;
        RECT 48.370 118.220 48.870 118.390 ;
        RECT 49.160 118.220 49.660 118.390 ;
        RECT 49.950 118.220 50.450 118.390 ;
        RECT 50.740 118.220 51.240 118.390 ;
        RECT 51.530 118.220 52.030 118.390 ;
        RECT 52.320 118.220 52.820 118.390 ;
        RECT 55.010 118.220 55.510 118.390 ;
        RECT 55.800 118.220 56.300 118.390 ;
        RECT 56.590 118.220 57.090 118.390 ;
        RECT 57.380 118.220 57.880 118.390 ;
        RECT 58.170 118.220 58.670 118.390 ;
        RECT 58.960 118.220 59.460 118.390 ;
        RECT 59.750 118.220 60.250 118.390 ;
        RECT 60.540 118.220 61.040 118.390 ;
        RECT 61.330 118.220 61.830 118.390 ;
        RECT 62.120 118.220 62.620 118.390 ;
        RECT 64.810 118.220 65.310 118.390 ;
        RECT 65.600 118.220 66.100 118.390 ;
        RECT 66.390 118.220 66.890 118.390 ;
        RECT 67.180 118.220 67.680 118.390 ;
        RECT 67.970 118.220 68.470 118.390 ;
        RECT 68.760 118.220 69.260 118.390 ;
        RECT 69.550 118.220 70.050 118.390 ;
        RECT 70.340 118.220 70.840 118.390 ;
        RECT 71.130 118.220 71.630 118.390 ;
        RECT 71.920 118.220 72.420 118.390 ;
        RECT 16.540 116.820 17.040 116.990 ;
        RECT 17.330 116.820 17.830 116.990 ;
        RECT 20.025 116.825 20.525 116.995 ;
        RECT 20.815 116.825 21.315 116.995 ;
        RECT 21.605 116.825 22.105 116.995 ;
        RECT 22.395 116.825 22.895 116.995 ;
        RECT 17.100 112.560 17.270 116.600 ;
        RECT 16.540 112.170 17.040 112.340 ;
        RECT 17.330 112.170 17.830 112.340 ;
        RECT 16.305 109.000 16.475 110.040 ;
        RECT 17.885 109.000 18.055 110.040 ;
        RECT 16.535 108.610 17.035 108.780 ;
        RECT 17.325 108.610 17.825 108.780 ;
        RECT 20.585 106.565 20.755 116.605 ;
        RECT 22.165 106.565 22.335 116.605 ;
        RECT 25.470 107.580 25.970 107.750 ;
        RECT 26.260 107.580 26.760 107.750 ;
        RECT 27.050 107.580 27.550 107.750 ;
        RECT 27.840 107.580 28.340 107.750 ;
        RECT 28.630 107.580 29.130 107.750 ;
        RECT 29.420 107.580 29.920 107.750 ;
        RECT 30.210 107.580 30.710 107.750 ;
        RECT 31.000 107.580 31.500 107.750 ;
        RECT 31.790 107.580 32.290 107.750 ;
        RECT 32.580 107.580 33.080 107.750 ;
        RECT 35.410 107.580 35.910 107.750 ;
        RECT 36.200 107.580 36.700 107.750 ;
        RECT 36.990 107.580 37.490 107.750 ;
        RECT 37.780 107.580 38.280 107.750 ;
        RECT 38.570 107.580 39.070 107.750 ;
        RECT 39.360 107.580 39.860 107.750 ;
        RECT 40.150 107.580 40.650 107.750 ;
        RECT 40.940 107.580 41.440 107.750 ;
        RECT 41.730 107.580 42.230 107.750 ;
        RECT 42.520 107.580 43.020 107.750 ;
        RECT 45.210 107.580 45.710 107.750 ;
        RECT 46.000 107.580 46.500 107.750 ;
        RECT 46.790 107.580 47.290 107.750 ;
        RECT 47.580 107.580 48.080 107.750 ;
        RECT 48.370 107.580 48.870 107.750 ;
        RECT 49.160 107.580 49.660 107.750 ;
        RECT 49.950 107.580 50.450 107.750 ;
        RECT 50.740 107.580 51.240 107.750 ;
        RECT 51.530 107.580 52.030 107.750 ;
        RECT 52.320 107.580 52.820 107.750 ;
        RECT 55.010 107.580 55.510 107.750 ;
        RECT 55.800 107.580 56.300 107.750 ;
        RECT 56.590 107.580 57.090 107.750 ;
        RECT 57.380 107.580 57.880 107.750 ;
        RECT 58.170 107.580 58.670 107.750 ;
        RECT 58.960 107.580 59.460 107.750 ;
        RECT 59.750 107.580 60.250 107.750 ;
        RECT 60.540 107.580 61.040 107.750 ;
        RECT 61.330 107.580 61.830 107.750 ;
        RECT 62.120 107.580 62.620 107.750 ;
        RECT 64.810 107.580 65.310 107.750 ;
        RECT 65.600 107.580 66.100 107.750 ;
        RECT 66.390 107.580 66.890 107.750 ;
        RECT 67.180 107.580 67.680 107.750 ;
        RECT 67.970 107.580 68.470 107.750 ;
        RECT 68.760 107.580 69.260 107.750 ;
        RECT 69.550 107.580 70.050 107.750 ;
        RECT 70.340 107.580 70.840 107.750 ;
        RECT 71.130 107.580 71.630 107.750 ;
        RECT 71.920 107.580 72.420 107.750 ;
        RECT 25.470 107.040 25.970 107.210 ;
        RECT 26.260 107.040 26.760 107.210 ;
        RECT 27.050 107.040 27.550 107.210 ;
        RECT 27.840 107.040 28.340 107.210 ;
        RECT 28.630 107.040 29.130 107.210 ;
        RECT 29.420 107.040 29.920 107.210 ;
        RECT 30.210 107.040 30.710 107.210 ;
        RECT 31.000 107.040 31.500 107.210 ;
        RECT 31.790 107.040 32.290 107.210 ;
        RECT 32.580 107.040 33.080 107.210 ;
        RECT 35.410 107.040 35.910 107.210 ;
        RECT 36.200 107.040 36.700 107.210 ;
        RECT 36.990 107.040 37.490 107.210 ;
        RECT 37.780 107.040 38.280 107.210 ;
        RECT 38.570 107.040 39.070 107.210 ;
        RECT 39.360 107.040 39.860 107.210 ;
        RECT 40.150 107.040 40.650 107.210 ;
        RECT 40.940 107.040 41.440 107.210 ;
        RECT 41.730 107.040 42.230 107.210 ;
        RECT 42.520 107.040 43.020 107.210 ;
        RECT 45.210 107.040 45.710 107.210 ;
        RECT 46.000 107.040 46.500 107.210 ;
        RECT 46.790 107.040 47.290 107.210 ;
        RECT 47.580 107.040 48.080 107.210 ;
        RECT 48.370 107.040 48.870 107.210 ;
        RECT 49.160 107.040 49.660 107.210 ;
        RECT 49.950 107.040 50.450 107.210 ;
        RECT 50.740 107.040 51.240 107.210 ;
        RECT 51.530 107.040 52.030 107.210 ;
        RECT 52.320 107.040 52.820 107.210 ;
        RECT 55.010 107.040 55.510 107.210 ;
        RECT 55.800 107.040 56.300 107.210 ;
        RECT 56.590 107.040 57.090 107.210 ;
        RECT 57.380 107.040 57.880 107.210 ;
        RECT 58.170 107.040 58.670 107.210 ;
        RECT 58.960 107.040 59.460 107.210 ;
        RECT 59.750 107.040 60.250 107.210 ;
        RECT 60.540 107.040 61.040 107.210 ;
        RECT 61.330 107.040 61.830 107.210 ;
        RECT 62.120 107.040 62.620 107.210 ;
        RECT 64.810 107.040 65.310 107.210 ;
        RECT 65.600 107.040 66.100 107.210 ;
        RECT 66.390 107.040 66.890 107.210 ;
        RECT 67.180 107.040 67.680 107.210 ;
        RECT 67.970 107.040 68.470 107.210 ;
        RECT 68.760 107.040 69.260 107.210 ;
        RECT 69.550 107.040 70.050 107.210 ;
        RECT 70.340 107.040 70.840 107.210 ;
        RECT 71.130 107.040 71.630 107.210 ;
        RECT 71.920 107.040 72.420 107.210 ;
        RECT 20.025 106.175 20.525 106.345 ;
        RECT 20.815 106.175 21.315 106.345 ;
        RECT 21.605 106.175 22.105 106.345 ;
        RECT 22.395 106.175 22.895 106.345 ;
        RECT 16.840 103.950 17.340 104.120 ;
        RECT 16.610 102.740 16.780 103.780 ;
        RECT 16.840 102.400 17.340 102.570 ;
        RECT 19.535 101.460 20.035 101.630 ;
        RECT 20.325 101.460 20.825 101.630 ;
        RECT 21.115 101.460 21.615 101.630 ;
        RECT 21.905 101.460 22.405 101.630 ;
        RECT 16.840 100.460 17.340 100.630 ;
        RECT 17.400 96.250 17.570 100.290 ;
        RECT 20.095 96.250 20.265 101.290 ;
        RECT 21.675 96.250 21.845 101.290 ;
        RECT 25.470 96.400 25.970 96.570 ;
        RECT 26.260 96.400 26.760 96.570 ;
        RECT 27.050 96.400 27.550 96.570 ;
        RECT 27.840 96.400 28.340 96.570 ;
        RECT 28.630 96.400 29.130 96.570 ;
        RECT 29.420 96.400 29.920 96.570 ;
        RECT 30.210 96.400 30.710 96.570 ;
        RECT 31.000 96.400 31.500 96.570 ;
        RECT 31.790 96.400 32.290 96.570 ;
        RECT 32.580 96.400 33.080 96.570 ;
        RECT 35.410 96.400 35.910 96.570 ;
        RECT 36.200 96.400 36.700 96.570 ;
        RECT 36.990 96.400 37.490 96.570 ;
        RECT 37.780 96.400 38.280 96.570 ;
        RECT 38.570 96.400 39.070 96.570 ;
        RECT 39.360 96.400 39.860 96.570 ;
        RECT 40.150 96.400 40.650 96.570 ;
        RECT 40.940 96.400 41.440 96.570 ;
        RECT 41.730 96.400 42.230 96.570 ;
        RECT 42.520 96.400 43.020 96.570 ;
        RECT 45.210 96.400 45.710 96.570 ;
        RECT 46.000 96.400 46.500 96.570 ;
        RECT 46.790 96.400 47.290 96.570 ;
        RECT 47.580 96.400 48.080 96.570 ;
        RECT 48.370 96.400 48.870 96.570 ;
        RECT 49.160 96.400 49.660 96.570 ;
        RECT 49.950 96.400 50.450 96.570 ;
        RECT 50.740 96.400 51.240 96.570 ;
        RECT 51.530 96.400 52.030 96.570 ;
        RECT 52.320 96.400 52.820 96.570 ;
        RECT 55.010 96.400 55.510 96.570 ;
        RECT 55.800 96.400 56.300 96.570 ;
        RECT 56.590 96.400 57.090 96.570 ;
        RECT 57.380 96.400 57.880 96.570 ;
        RECT 58.170 96.400 58.670 96.570 ;
        RECT 58.960 96.400 59.460 96.570 ;
        RECT 59.750 96.400 60.250 96.570 ;
        RECT 60.540 96.400 61.040 96.570 ;
        RECT 61.330 96.400 61.830 96.570 ;
        RECT 62.120 96.400 62.620 96.570 ;
        RECT 64.810 96.400 65.310 96.570 ;
        RECT 65.600 96.400 66.100 96.570 ;
        RECT 66.390 96.400 66.890 96.570 ;
        RECT 67.180 96.400 67.680 96.570 ;
        RECT 67.970 96.400 68.470 96.570 ;
        RECT 68.760 96.400 69.260 96.570 ;
        RECT 69.550 96.400 70.050 96.570 ;
        RECT 70.340 96.400 70.840 96.570 ;
        RECT 71.130 96.400 71.630 96.570 ;
        RECT 71.920 96.400 72.420 96.570 ;
        RECT 16.840 95.910 17.340 96.080 ;
        RECT 19.535 95.910 20.035 96.080 ;
        RECT 20.325 95.910 20.825 96.080 ;
        RECT 21.115 95.910 21.615 96.080 ;
        RECT 21.905 95.910 22.405 96.080 ;
        RECT 15.285 93.950 15.785 94.120 ;
        RECT 16.075 93.950 16.575 94.120 ;
        RECT 16.865 93.950 17.365 94.120 ;
        RECT 17.655 93.950 18.155 94.120 ;
        RECT 18.445 93.950 18.945 94.120 ;
        RECT 19.235 93.950 19.735 94.120 ;
        RECT 20.025 93.950 20.525 94.120 ;
        RECT 20.815 93.950 21.315 94.120 ;
        RECT 21.605 93.950 22.105 94.120 ;
        RECT 22.395 93.950 22.895 94.120 ;
        RECT 25.475 93.965 25.975 94.135 ;
        RECT 26.265 93.965 26.765 94.135 ;
        RECT 27.055 93.965 27.555 94.135 ;
        RECT 27.845 93.965 28.345 94.135 ;
        RECT 28.635 93.965 29.135 94.135 ;
        RECT 29.425 93.965 29.925 94.135 ;
        RECT 30.215 93.965 30.715 94.135 ;
        RECT 31.005 93.965 31.505 94.135 ;
        RECT 31.795 93.965 32.295 94.135 ;
        RECT 32.585 93.965 33.085 94.135 ;
        RECT 35.415 93.965 35.915 94.135 ;
        RECT 36.205 93.965 36.705 94.135 ;
        RECT 36.995 93.965 37.495 94.135 ;
        RECT 37.785 93.965 38.285 94.135 ;
        RECT 38.575 93.965 39.075 94.135 ;
        RECT 39.365 93.965 39.865 94.135 ;
        RECT 40.155 93.965 40.655 94.135 ;
        RECT 40.945 93.965 41.445 94.135 ;
        RECT 41.735 93.965 42.235 94.135 ;
        RECT 42.525 93.965 43.025 94.135 ;
        RECT 45.215 93.965 45.715 94.135 ;
        RECT 46.005 93.965 46.505 94.135 ;
        RECT 46.795 93.965 47.295 94.135 ;
        RECT 47.585 93.965 48.085 94.135 ;
        RECT 48.375 93.965 48.875 94.135 ;
        RECT 49.165 93.965 49.665 94.135 ;
        RECT 49.955 93.965 50.455 94.135 ;
        RECT 50.745 93.965 51.245 94.135 ;
        RECT 51.535 93.965 52.035 94.135 ;
        RECT 52.325 93.965 52.825 94.135 ;
        RECT 55.015 93.965 55.515 94.135 ;
        RECT 55.805 93.965 56.305 94.135 ;
        RECT 56.595 93.965 57.095 94.135 ;
        RECT 57.385 93.965 57.885 94.135 ;
        RECT 58.175 93.965 58.675 94.135 ;
        RECT 58.965 93.965 59.465 94.135 ;
        RECT 59.755 93.965 60.255 94.135 ;
        RECT 60.545 93.965 61.045 94.135 ;
        RECT 61.335 93.965 61.835 94.135 ;
        RECT 62.125 93.965 62.625 94.135 ;
        RECT 64.815 93.965 65.315 94.135 ;
        RECT 65.605 93.965 66.105 94.135 ;
        RECT 66.395 93.965 66.895 94.135 ;
        RECT 67.185 93.965 67.685 94.135 ;
        RECT 67.975 93.965 68.475 94.135 ;
        RECT 68.765 93.965 69.265 94.135 ;
        RECT 69.555 93.965 70.055 94.135 ;
        RECT 70.345 93.965 70.845 94.135 ;
        RECT 71.135 93.965 71.635 94.135 ;
        RECT 71.925 93.965 72.425 94.135 ;
        RECT 15.845 83.740 16.015 93.780 ;
        RECT 17.425 83.740 17.595 93.780 ;
        RECT 19.005 83.740 19.175 93.780 ;
        RECT 20.585 83.740 20.755 93.780 ;
        RECT 22.165 83.740 22.335 93.780 ;
        RECT 15.285 83.400 15.785 83.570 ;
        RECT 16.075 83.400 16.575 83.570 ;
        RECT 16.865 83.400 17.365 83.570 ;
        RECT 17.655 83.400 18.155 83.570 ;
        RECT 18.445 83.400 18.945 83.570 ;
        RECT 19.235 83.400 19.735 83.570 ;
        RECT 20.025 83.400 20.525 83.570 ;
        RECT 20.815 83.400 21.315 83.570 ;
        RECT 21.605 83.400 22.105 83.570 ;
        RECT 22.395 83.400 22.895 83.570 ;
        RECT 25.475 83.415 25.975 83.585 ;
        RECT 26.265 83.415 26.765 83.585 ;
        RECT 27.055 83.415 27.555 83.585 ;
        RECT 27.845 83.415 28.345 83.585 ;
        RECT 28.635 83.415 29.135 83.585 ;
        RECT 29.425 83.415 29.925 83.585 ;
        RECT 30.215 83.415 30.715 83.585 ;
        RECT 31.005 83.415 31.505 83.585 ;
        RECT 31.795 83.415 32.295 83.585 ;
        RECT 32.585 83.415 33.085 83.585 ;
        RECT 35.415 83.415 35.915 83.585 ;
        RECT 36.205 83.415 36.705 83.585 ;
        RECT 36.995 83.415 37.495 83.585 ;
        RECT 37.785 83.415 38.285 83.585 ;
        RECT 38.575 83.415 39.075 83.585 ;
        RECT 39.365 83.415 39.865 83.585 ;
        RECT 40.155 83.415 40.655 83.585 ;
        RECT 40.945 83.415 41.445 83.585 ;
        RECT 41.735 83.415 42.235 83.585 ;
        RECT 42.525 83.415 43.025 83.585 ;
        RECT 45.215 83.415 45.715 83.585 ;
        RECT 46.005 83.415 46.505 83.585 ;
        RECT 46.795 83.415 47.295 83.585 ;
        RECT 47.585 83.415 48.085 83.585 ;
        RECT 48.375 83.415 48.875 83.585 ;
        RECT 49.165 83.415 49.665 83.585 ;
        RECT 49.955 83.415 50.455 83.585 ;
        RECT 50.745 83.415 51.245 83.585 ;
        RECT 51.535 83.415 52.035 83.585 ;
        RECT 52.325 83.415 52.825 83.585 ;
        RECT 55.015 83.415 55.515 83.585 ;
        RECT 55.805 83.415 56.305 83.585 ;
        RECT 56.595 83.415 57.095 83.585 ;
        RECT 57.385 83.415 57.885 83.585 ;
        RECT 58.175 83.415 58.675 83.585 ;
        RECT 58.965 83.415 59.465 83.585 ;
        RECT 59.755 83.415 60.255 83.585 ;
        RECT 60.545 83.415 61.045 83.585 ;
        RECT 61.335 83.415 61.835 83.585 ;
        RECT 62.125 83.415 62.625 83.585 ;
        RECT 64.815 83.415 65.315 83.585 ;
        RECT 65.605 83.415 66.105 83.585 ;
        RECT 66.395 83.415 66.895 83.585 ;
        RECT 67.185 83.415 67.685 83.585 ;
        RECT 67.975 83.415 68.475 83.585 ;
        RECT 68.765 83.415 69.265 83.585 ;
        RECT 69.555 83.415 70.055 83.585 ;
        RECT 70.345 83.415 70.845 83.585 ;
        RECT 71.135 83.415 71.635 83.585 ;
        RECT 71.925 83.415 72.425 83.585 ;
        RECT 25.475 82.885 25.975 83.055 ;
        RECT 26.265 82.885 26.765 83.055 ;
        RECT 27.055 82.885 27.555 83.055 ;
        RECT 27.845 82.885 28.345 83.055 ;
        RECT 28.635 82.885 29.135 83.055 ;
        RECT 29.425 82.885 29.925 83.055 ;
        RECT 30.215 82.885 30.715 83.055 ;
        RECT 31.005 82.885 31.505 83.055 ;
        RECT 31.795 82.885 32.295 83.055 ;
        RECT 32.585 82.885 33.085 83.055 ;
        RECT 35.415 82.885 35.915 83.055 ;
        RECT 36.205 82.885 36.705 83.055 ;
        RECT 36.995 82.885 37.495 83.055 ;
        RECT 37.785 82.885 38.285 83.055 ;
        RECT 38.575 82.885 39.075 83.055 ;
        RECT 39.365 82.885 39.865 83.055 ;
        RECT 40.155 82.885 40.655 83.055 ;
        RECT 40.945 82.885 41.445 83.055 ;
        RECT 41.735 82.885 42.235 83.055 ;
        RECT 42.525 82.885 43.025 83.055 ;
        RECT 45.215 82.885 45.715 83.055 ;
        RECT 46.005 82.885 46.505 83.055 ;
        RECT 46.795 82.885 47.295 83.055 ;
        RECT 47.585 82.885 48.085 83.055 ;
        RECT 48.375 82.885 48.875 83.055 ;
        RECT 49.165 82.885 49.665 83.055 ;
        RECT 49.955 82.885 50.455 83.055 ;
        RECT 50.745 82.885 51.245 83.055 ;
        RECT 51.535 82.885 52.035 83.055 ;
        RECT 52.325 82.885 52.825 83.055 ;
        RECT 55.015 82.885 55.515 83.055 ;
        RECT 55.805 82.885 56.305 83.055 ;
        RECT 56.595 82.885 57.095 83.055 ;
        RECT 57.385 82.885 57.885 83.055 ;
        RECT 58.175 82.885 58.675 83.055 ;
        RECT 58.965 82.885 59.465 83.055 ;
        RECT 59.755 82.885 60.255 83.055 ;
        RECT 60.545 82.885 61.045 83.055 ;
        RECT 61.335 82.885 61.835 83.055 ;
        RECT 62.125 82.885 62.625 83.055 ;
        RECT 64.815 82.885 65.315 83.055 ;
        RECT 65.605 82.885 66.105 83.055 ;
        RECT 66.395 82.885 66.895 83.055 ;
        RECT 67.185 82.885 67.685 83.055 ;
        RECT 67.975 82.885 68.475 83.055 ;
        RECT 68.765 82.885 69.265 83.055 ;
        RECT 69.555 82.885 70.055 83.055 ;
        RECT 70.345 82.885 70.845 83.055 ;
        RECT 71.135 82.885 71.635 83.055 ;
        RECT 71.925 82.885 72.425 83.055 ;
        RECT 3.595 80.690 4.095 80.860 ;
        RECT 4.385 80.690 4.885 80.860 ;
        RECT 5.175 80.690 5.675 80.860 ;
        RECT 5.965 80.690 6.465 80.860 ;
        RECT 6.755 80.690 7.255 80.860 ;
        RECT 8.885 80.690 9.385 80.860 ;
        RECT 9.675 80.690 10.175 80.860 ;
        RECT 10.465 80.690 10.965 80.860 ;
        RECT 11.255 80.690 11.755 80.860 ;
        RECT 12.045 80.690 12.545 80.860 ;
        RECT 4.155 78.430 4.325 80.470 ;
        RECT 5.735 78.430 5.905 80.470 ;
        RECT 7.315 78.430 7.485 80.470 ;
        RECT 8.655 78.430 8.825 80.470 ;
        RECT 10.235 78.430 10.405 80.470 ;
        RECT 11.815 78.430 11.985 80.470 ;
        RECT 17.965 80.110 18.465 80.280 ;
        RECT 18.755 80.110 19.255 80.280 ;
        RECT 21.045 80.110 21.545 80.280 ;
        RECT 21.835 80.110 22.335 80.280 ;
        RECT 3.595 78.040 4.095 78.210 ;
        RECT 4.385 78.040 4.885 78.210 ;
        RECT 5.175 78.040 5.675 78.210 ;
        RECT 5.965 78.040 6.465 78.210 ;
        RECT 6.755 78.040 7.255 78.210 ;
        RECT 8.885 78.040 9.385 78.210 ;
        RECT 9.675 78.040 10.175 78.210 ;
        RECT 10.465 78.040 10.965 78.210 ;
        RECT 11.255 78.040 11.755 78.210 ;
        RECT 12.045 78.040 12.545 78.210 ;
        RECT 1.015 65.295 1.185 75.335 ;
        RECT 2.205 65.295 2.375 75.335 ;
        RECT 3.395 65.295 3.565 75.335 ;
        RECT 4.585 65.295 4.755 75.335 ;
        RECT 5.775 65.295 5.945 75.335 ;
        RECT 6.965 65.295 7.135 75.335 ;
        RECT 8.865 65.295 9.035 75.335 ;
        RECT 10.055 65.295 10.225 75.335 ;
        RECT 11.245 65.295 11.415 75.335 ;
        RECT 12.435 65.295 12.605 75.335 ;
        RECT 13.625 65.295 13.795 75.335 ;
        RECT 14.815 65.295 14.985 75.335 ;
        RECT 18.525 69.850 18.695 79.890 ;
        RECT 21.605 69.850 21.775 79.890 ;
        RECT 25.475 72.335 25.975 72.505 ;
        RECT 26.265 72.335 26.765 72.505 ;
        RECT 27.055 72.335 27.555 72.505 ;
        RECT 27.845 72.335 28.345 72.505 ;
        RECT 28.635 72.335 29.135 72.505 ;
        RECT 29.425 72.335 29.925 72.505 ;
        RECT 30.215 72.335 30.715 72.505 ;
        RECT 31.005 72.335 31.505 72.505 ;
        RECT 31.795 72.335 32.295 72.505 ;
        RECT 32.585 72.335 33.085 72.505 ;
        RECT 35.415 72.335 35.915 72.505 ;
        RECT 36.205 72.335 36.705 72.505 ;
        RECT 36.995 72.335 37.495 72.505 ;
        RECT 37.785 72.335 38.285 72.505 ;
        RECT 38.575 72.335 39.075 72.505 ;
        RECT 39.365 72.335 39.865 72.505 ;
        RECT 40.155 72.335 40.655 72.505 ;
        RECT 40.945 72.335 41.445 72.505 ;
        RECT 41.735 72.335 42.235 72.505 ;
        RECT 42.525 72.335 43.025 72.505 ;
        RECT 45.215 72.335 45.715 72.505 ;
        RECT 46.005 72.335 46.505 72.505 ;
        RECT 46.795 72.335 47.295 72.505 ;
        RECT 47.585 72.335 48.085 72.505 ;
        RECT 48.375 72.335 48.875 72.505 ;
        RECT 49.165 72.335 49.665 72.505 ;
        RECT 49.955 72.335 50.455 72.505 ;
        RECT 50.745 72.335 51.245 72.505 ;
        RECT 51.535 72.335 52.035 72.505 ;
        RECT 52.325 72.335 52.825 72.505 ;
        RECT 55.015 72.335 55.515 72.505 ;
        RECT 55.805 72.335 56.305 72.505 ;
        RECT 56.595 72.335 57.095 72.505 ;
        RECT 57.385 72.335 57.885 72.505 ;
        RECT 58.175 72.335 58.675 72.505 ;
        RECT 58.965 72.335 59.465 72.505 ;
        RECT 59.755 72.335 60.255 72.505 ;
        RECT 60.545 72.335 61.045 72.505 ;
        RECT 61.335 72.335 61.835 72.505 ;
        RECT 62.125 72.335 62.625 72.505 ;
        RECT 64.815 72.335 65.315 72.505 ;
        RECT 65.605 72.335 66.105 72.505 ;
        RECT 66.395 72.335 66.895 72.505 ;
        RECT 67.185 72.335 67.685 72.505 ;
        RECT 67.975 72.335 68.475 72.505 ;
        RECT 68.765 72.335 69.265 72.505 ;
        RECT 69.555 72.335 70.055 72.505 ;
        RECT 70.345 72.335 70.845 72.505 ;
        RECT 71.135 72.335 71.635 72.505 ;
        RECT 71.925 72.335 72.425 72.505 ;
        RECT 17.965 69.460 18.465 69.630 ;
        RECT 18.755 69.460 19.255 69.630 ;
        RECT 21.045 69.460 21.545 69.630 ;
        RECT 21.835 69.460 22.335 69.630 ;
        RECT 25.475 69.325 25.975 69.495 ;
        RECT 26.265 69.325 26.765 69.495 ;
        RECT 27.055 69.325 27.555 69.495 ;
        RECT 27.845 69.325 28.345 69.495 ;
        RECT 28.635 69.325 29.135 69.495 ;
        RECT 29.425 69.325 29.925 69.495 ;
        RECT 30.215 69.325 30.715 69.495 ;
        RECT 31.005 69.325 31.505 69.495 ;
        RECT 31.795 69.325 32.295 69.495 ;
        RECT 32.585 69.325 33.085 69.495 ;
        RECT 35.415 69.325 35.915 69.495 ;
        RECT 36.205 69.325 36.705 69.495 ;
        RECT 36.995 69.325 37.495 69.495 ;
        RECT 37.785 69.325 38.285 69.495 ;
        RECT 38.575 69.325 39.075 69.495 ;
        RECT 39.365 69.325 39.865 69.495 ;
        RECT 40.155 69.325 40.655 69.495 ;
        RECT 40.945 69.325 41.445 69.495 ;
        RECT 41.735 69.325 42.235 69.495 ;
        RECT 42.525 69.325 43.025 69.495 ;
        RECT 45.215 69.325 45.715 69.495 ;
        RECT 46.005 69.325 46.505 69.495 ;
        RECT 46.795 69.325 47.295 69.495 ;
        RECT 47.585 69.325 48.085 69.495 ;
        RECT 48.375 69.325 48.875 69.495 ;
        RECT 49.165 69.325 49.665 69.495 ;
        RECT 49.955 69.325 50.455 69.495 ;
        RECT 50.745 69.325 51.245 69.495 ;
        RECT 51.535 69.325 52.035 69.495 ;
        RECT 52.325 69.325 52.825 69.495 ;
        RECT 55.015 69.325 55.515 69.495 ;
        RECT 55.805 69.325 56.305 69.495 ;
        RECT 56.595 69.325 57.095 69.495 ;
        RECT 57.385 69.325 57.885 69.495 ;
        RECT 58.175 69.325 58.675 69.495 ;
        RECT 58.965 69.325 59.465 69.495 ;
        RECT 59.755 69.325 60.255 69.495 ;
        RECT 60.545 69.325 61.045 69.495 ;
        RECT 61.335 69.325 61.835 69.495 ;
        RECT 62.125 69.325 62.625 69.495 ;
        RECT 64.815 69.325 65.315 69.495 ;
        RECT 65.605 69.325 66.105 69.495 ;
        RECT 66.395 69.325 66.895 69.495 ;
        RECT 67.185 69.325 67.685 69.495 ;
        RECT 67.975 69.325 68.475 69.495 ;
        RECT 68.765 69.325 69.265 69.495 ;
        RECT 69.555 69.325 70.055 69.495 ;
        RECT 70.345 69.325 70.845 69.495 ;
        RECT 71.135 69.325 71.635 69.495 ;
        RECT 71.925 69.325 72.425 69.495 ;
        RECT 17.965 67.030 18.465 67.200 ;
        RECT 18.755 67.030 19.255 67.200 ;
        RECT 21.045 67.030 21.545 67.200 ;
        RECT 21.835 67.030 22.335 67.200 ;
        RECT 3.105 60.730 3.275 62.770 ;
        RECT 4.065 60.730 4.235 62.770 ;
        RECT 5.025 60.730 5.195 62.770 ;
        RECT 5.975 60.730 6.145 62.770 ;
        RECT 6.935 60.730 7.105 62.770 ;
        RECT 9.035 60.730 9.205 62.770 ;
        RECT 9.995 60.730 10.165 62.770 ;
        RECT 10.955 60.730 11.125 62.770 ;
        RECT 11.905 60.730 12.075 62.770 ;
        RECT 12.865 60.730 13.035 62.770 ;
        RECT 18.525 61.820 18.695 66.860 ;
        RECT 21.605 61.820 21.775 66.860 ;
        RECT 17.965 61.480 18.465 61.650 ;
        RECT 18.755 61.480 19.255 61.650 ;
        RECT 21.045 61.480 21.545 61.650 ;
        RECT 21.835 61.480 22.335 61.650 ;
        RECT 25.475 58.775 25.975 58.945 ;
        RECT 26.265 58.775 26.765 58.945 ;
        RECT 27.055 58.775 27.555 58.945 ;
        RECT 27.845 58.775 28.345 58.945 ;
        RECT 28.635 58.775 29.135 58.945 ;
        RECT 29.425 58.775 29.925 58.945 ;
        RECT 30.215 58.775 30.715 58.945 ;
        RECT 31.005 58.775 31.505 58.945 ;
        RECT 31.795 58.775 32.295 58.945 ;
        RECT 32.585 58.775 33.085 58.945 ;
        RECT 35.415 58.775 35.915 58.945 ;
        RECT 36.205 58.775 36.705 58.945 ;
        RECT 36.995 58.775 37.495 58.945 ;
        RECT 37.785 58.775 38.285 58.945 ;
        RECT 38.575 58.775 39.075 58.945 ;
        RECT 39.365 58.775 39.865 58.945 ;
        RECT 40.155 58.775 40.655 58.945 ;
        RECT 40.945 58.775 41.445 58.945 ;
        RECT 41.735 58.775 42.235 58.945 ;
        RECT 42.525 58.775 43.025 58.945 ;
        RECT 45.215 58.775 45.715 58.945 ;
        RECT 46.005 58.775 46.505 58.945 ;
        RECT 46.795 58.775 47.295 58.945 ;
        RECT 47.585 58.775 48.085 58.945 ;
        RECT 48.375 58.775 48.875 58.945 ;
        RECT 49.165 58.775 49.665 58.945 ;
        RECT 49.955 58.775 50.455 58.945 ;
        RECT 50.745 58.775 51.245 58.945 ;
        RECT 51.535 58.775 52.035 58.945 ;
        RECT 52.325 58.775 52.825 58.945 ;
        RECT 55.015 58.775 55.515 58.945 ;
        RECT 55.805 58.775 56.305 58.945 ;
        RECT 56.595 58.775 57.095 58.945 ;
        RECT 57.385 58.775 57.885 58.945 ;
        RECT 58.175 58.775 58.675 58.945 ;
        RECT 58.965 58.775 59.465 58.945 ;
        RECT 59.755 58.775 60.255 58.945 ;
        RECT 60.545 58.775 61.045 58.945 ;
        RECT 61.335 58.775 61.835 58.945 ;
        RECT 62.125 58.775 62.625 58.945 ;
        RECT 64.815 58.775 65.315 58.945 ;
        RECT 65.605 58.775 66.105 58.945 ;
        RECT 66.395 58.775 66.895 58.945 ;
        RECT 67.185 58.775 67.685 58.945 ;
        RECT 67.975 58.775 68.475 58.945 ;
        RECT 68.765 58.775 69.265 58.945 ;
        RECT 69.555 58.775 70.055 58.945 ;
        RECT 70.345 58.775 70.845 58.945 ;
        RECT 71.135 58.775 71.635 58.945 ;
        RECT 71.925 58.775 72.425 58.945 ;
        RECT 15.285 58.260 15.785 58.430 ;
        RECT 16.075 58.260 16.575 58.430 ;
        RECT 16.865 58.260 17.365 58.430 ;
        RECT 17.655 58.260 18.155 58.430 ;
        RECT 18.445 58.260 18.945 58.430 ;
        RECT 19.235 58.260 19.735 58.430 ;
        RECT 20.025 58.260 20.525 58.430 ;
        RECT 20.815 58.260 21.315 58.430 ;
        RECT 21.605 58.260 22.105 58.430 ;
        RECT 22.395 58.260 22.895 58.430 ;
        RECT 25.475 58.245 25.975 58.415 ;
        RECT 26.265 58.245 26.765 58.415 ;
        RECT 27.055 58.245 27.555 58.415 ;
        RECT 27.845 58.245 28.345 58.415 ;
        RECT 28.635 58.245 29.135 58.415 ;
        RECT 29.425 58.245 29.925 58.415 ;
        RECT 30.215 58.245 30.715 58.415 ;
        RECT 31.005 58.245 31.505 58.415 ;
        RECT 31.795 58.245 32.295 58.415 ;
        RECT 32.585 58.245 33.085 58.415 ;
        RECT 35.415 58.245 35.915 58.415 ;
        RECT 36.205 58.245 36.705 58.415 ;
        RECT 36.995 58.245 37.495 58.415 ;
        RECT 37.785 58.245 38.285 58.415 ;
        RECT 38.575 58.245 39.075 58.415 ;
        RECT 39.365 58.245 39.865 58.415 ;
        RECT 40.155 58.245 40.655 58.415 ;
        RECT 40.945 58.245 41.445 58.415 ;
        RECT 41.735 58.245 42.235 58.415 ;
        RECT 42.525 58.245 43.025 58.415 ;
        RECT 45.215 58.245 45.715 58.415 ;
        RECT 46.005 58.245 46.505 58.415 ;
        RECT 46.795 58.245 47.295 58.415 ;
        RECT 47.585 58.245 48.085 58.415 ;
        RECT 48.375 58.245 48.875 58.415 ;
        RECT 49.165 58.245 49.665 58.415 ;
        RECT 49.955 58.245 50.455 58.415 ;
        RECT 50.745 58.245 51.245 58.415 ;
        RECT 51.535 58.245 52.035 58.415 ;
        RECT 52.325 58.245 52.825 58.415 ;
        RECT 55.015 58.245 55.515 58.415 ;
        RECT 55.805 58.245 56.305 58.415 ;
        RECT 56.595 58.245 57.095 58.415 ;
        RECT 57.385 58.245 57.885 58.415 ;
        RECT 58.175 58.245 58.675 58.415 ;
        RECT 58.965 58.245 59.465 58.415 ;
        RECT 59.755 58.245 60.255 58.415 ;
        RECT 60.545 58.245 61.045 58.415 ;
        RECT 61.335 58.245 61.835 58.415 ;
        RECT 62.125 58.245 62.625 58.415 ;
        RECT 64.815 58.245 65.315 58.415 ;
        RECT 65.605 58.245 66.105 58.415 ;
        RECT 66.395 58.245 66.895 58.415 ;
        RECT 67.185 58.245 67.685 58.415 ;
        RECT 67.975 58.245 68.475 58.415 ;
        RECT 68.765 58.245 69.265 58.415 ;
        RECT 69.555 58.245 70.055 58.415 ;
        RECT 70.345 58.245 70.845 58.415 ;
        RECT 71.135 58.245 71.635 58.415 ;
        RECT 71.925 58.245 72.425 58.415 ;
        RECT 15.845 48.050 16.015 58.090 ;
        RECT 17.425 48.050 17.595 58.090 ;
        RECT 19.005 48.050 19.175 58.090 ;
        RECT 20.585 48.050 20.755 58.090 ;
        RECT 22.165 48.050 22.335 58.090 ;
        RECT 15.285 47.710 15.785 47.880 ;
        RECT 16.075 47.710 16.575 47.880 ;
        RECT 16.865 47.710 17.365 47.880 ;
        RECT 17.655 47.710 18.155 47.880 ;
        RECT 18.445 47.710 18.945 47.880 ;
        RECT 19.235 47.710 19.735 47.880 ;
        RECT 20.025 47.710 20.525 47.880 ;
        RECT 20.815 47.710 21.315 47.880 ;
        RECT 21.605 47.710 22.105 47.880 ;
        RECT 22.395 47.710 22.895 47.880 ;
        RECT 25.475 47.695 25.975 47.865 ;
        RECT 26.265 47.695 26.765 47.865 ;
        RECT 27.055 47.695 27.555 47.865 ;
        RECT 27.845 47.695 28.345 47.865 ;
        RECT 28.635 47.695 29.135 47.865 ;
        RECT 29.425 47.695 29.925 47.865 ;
        RECT 30.215 47.695 30.715 47.865 ;
        RECT 31.005 47.695 31.505 47.865 ;
        RECT 31.795 47.695 32.295 47.865 ;
        RECT 32.585 47.695 33.085 47.865 ;
        RECT 35.415 47.695 35.915 47.865 ;
        RECT 36.205 47.695 36.705 47.865 ;
        RECT 36.995 47.695 37.495 47.865 ;
        RECT 37.785 47.695 38.285 47.865 ;
        RECT 38.575 47.695 39.075 47.865 ;
        RECT 39.365 47.695 39.865 47.865 ;
        RECT 40.155 47.695 40.655 47.865 ;
        RECT 40.945 47.695 41.445 47.865 ;
        RECT 41.735 47.695 42.235 47.865 ;
        RECT 42.525 47.695 43.025 47.865 ;
        RECT 45.215 47.695 45.715 47.865 ;
        RECT 46.005 47.695 46.505 47.865 ;
        RECT 46.795 47.695 47.295 47.865 ;
        RECT 47.585 47.695 48.085 47.865 ;
        RECT 48.375 47.695 48.875 47.865 ;
        RECT 49.165 47.695 49.665 47.865 ;
        RECT 49.955 47.695 50.455 47.865 ;
        RECT 50.745 47.695 51.245 47.865 ;
        RECT 51.535 47.695 52.035 47.865 ;
        RECT 52.325 47.695 52.825 47.865 ;
        RECT 55.015 47.695 55.515 47.865 ;
        RECT 55.805 47.695 56.305 47.865 ;
        RECT 56.595 47.695 57.095 47.865 ;
        RECT 57.385 47.695 57.885 47.865 ;
        RECT 58.175 47.695 58.675 47.865 ;
        RECT 58.965 47.695 59.465 47.865 ;
        RECT 59.755 47.695 60.255 47.865 ;
        RECT 60.545 47.695 61.045 47.865 ;
        RECT 61.335 47.695 61.835 47.865 ;
        RECT 62.125 47.695 62.625 47.865 ;
        RECT 64.815 47.695 65.315 47.865 ;
        RECT 65.605 47.695 66.105 47.865 ;
        RECT 66.395 47.695 66.895 47.865 ;
        RECT 67.185 47.695 67.685 47.865 ;
        RECT 67.975 47.695 68.475 47.865 ;
        RECT 68.765 47.695 69.265 47.865 ;
        RECT 69.555 47.695 70.055 47.865 ;
        RECT 70.345 47.695 70.845 47.865 ;
        RECT 71.135 47.695 71.635 47.865 ;
        RECT 71.925 47.695 72.425 47.865 ;
        RECT 16.840 45.750 17.340 45.920 ;
        RECT 19.535 45.750 20.035 45.920 ;
        RECT 20.325 45.750 20.825 45.920 ;
        RECT 21.115 45.750 21.615 45.920 ;
        RECT 21.905 45.750 22.405 45.920 ;
        RECT 17.400 41.540 17.570 45.580 ;
        RECT 16.840 41.200 17.340 41.370 ;
        RECT 20.095 40.540 20.265 45.580 ;
        RECT 21.675 40.540 21.845 45.580 ;
        RECT 25.470 45.260 25.970 45.430 ;
        RECT 26.260 45.260 26.760 45.430 ;
        RECT 27.050 45.260 27.550 45.430 ;
        RECT 27.840 45.260 28.340 45.430 ;
        RECT 28.630 45.260 29.130 45.430 ;
        RECT 29.420 45.260 29.920 45.430 ;
        RECT 30.210 45.260 30.710 45.430 ;
        RECT 31.000 45.260 31.500 45.430 ;
        RECT 31.790 45.260 32.290 45.430 ;
        RECT 32.580 45.260 33.080 45.430 ;
        RECT 35.410 45.260 35.910 45.430 ;
        RECT 36.200 45.260 36.700 45.430 ;
        RECT 36.990 45.260 37.490 45.430 ;
        RECT 37.780 45.260 38.280 45.430 ;
        RECT 38.570 45.260 39.070 45.430 ;
        RECT 39.360 45.260 39.860 45.430 ;
        RECT 40.150 45.260 40.650 45.430 ;
        RECT 40.940 45.260 41.440 45.430 ;
        RECT 41.730 45.260 42.230 45.430 ;
        RECT 42.520 45.260 43.020 45.430 ;
        RECT 45.210 45.260 45.710 45.430 ;
        RECT 46.000 45.260 46.500 45.430 ;
        RECT 46.790 45.260 47.290 45.430 ;
        RECT 47.580 45.260 48.080 45.430 ;
        RECT 48.370 45.260 48.870 45.430 ;
        RECT 49.160 45.260 49.660 45.430 ;
        RECT 49.950 45.260 50.450 45.430 ;
        RECT 50.740 45.260 51.240 45.430 ;
        RECT 51.530 45.260 52.030 45.430 ;
        RECT 52.320 45.260 52.820 45.430 ;
        RECT 55.010 45.260 55.510 45.430 ;
        RECT 55.800 45.260 56.300 45.430 ;
        RECT 56.590 45.260 57.090 45.430 ;
        RECT 57.380 45.260 57.880 45.430 ;
        RECT 58.170 45.260 58.670 45.430 ;
        RECT 58.960 45.260 59.460 45.430 ;
        RECT 59.750 45.260 60.250 45.430 ;
        RECT 60.540 45.260 61.040 45.430 ;
        RECT 61.330 45.260 61.830 45.430 ;
        RECT 62.120 45.260 62.620 45.430 ;
        RECT 64.810 45.260 65.310 45.430 ;
        RECT 65.600 45.260 66.100 45.430 ;
        RECT 66.390 45.260 66.890 45.430 ;
        RECT 67.180 45.260 67.680 45.430 ;
        RECT 67.970 45.260 68.470 45.430 ;
        RECT 68.760 45.260 69.260 45.430 ;
        RECT 69.550 45.260 70.050 45.430 ;
        RECT 70.340 45.260 70.840 45.430 ;
        RECT 71.130 45.260 71.630 45.430 ;
        RECT 71.920 45.260 72.420 45.430 ;
        RECT 19.535 40.200 20.035 40.370 ;
        RECT 20.325 40.200 20.825 40.370 ;
        RECT 21.115 40.200 21.615 40.370 ;
        RECT 21.905 40.200 22.405 40.370 ;
        RECT 16.840 39.260 17.340 39.430 ;
        RECT 16.610 38.050 16.780 39.090 ;
        RECT 16.840 37.710 17.340 37.880 ;
        RECT 20.025 35.485 20.525 35.655 ;
        RECT 20.815 35.485 21.315 35.655 ;
        RECT 21.605 35.485 22.105 35.655 ;
        RECT 22.395 35.485 22.895 35.655 ;
        RECT 16.535 33.050 17.035 33.220 ;
        RECT 17.325 33.050 17.825 33.220 ;
        RECT 16.305 31.790 16.475 32.830 ;
        RECT 17.885 31.790 18.055 32.830 ;
        RECT 16.540 29.490 17.040 29.660 ;
        RECT 17.330 29.490 17.830 29.660 ;
        RECT 17.100 25.230 17.270 29.270 ;
        RECT 20.585 25.225 20.755 35.265 ;
        RECT 22.165 25.225 22.335 35.265 ;
        RECT 25.470 34.620 25.970 34.790 ;
        RECT 26.260 34.620 26.760 34.790 ;
        RECT 27.050 34.620 27.550 34.790 ;
        RECT 27.840 34.620 28.340 34.790 ;
        RECT 28.630 34.620 29.130 34.790 ;
        RECT 29.420 34.620 29.920 34.790 ;
        RECT 30.210 34.620 30.710 34.790 ;
        RECT 31.000 34.620 31.500 34.790 ;
        RECT 31.790 34.620 32.290 34.790 ;
        RECT 32.580 34.620 33.080 34.790 ;
        RECT 35.410 34.620 35.910 34.790 ;
        RECT 36.200 34.620 36.700 34.790 ;
        RECT 36.990 34.620 37.490 34.790 ;
        RECT 37.780 34.620 38.280 34.790 ;
        RECT 38.570 34.620 39.070 34.790 ;
        RECT 39.360 34.620 39.860 34.790 ;
        RECT 40.150 34.620 40.650 34.790 ;
        RECT 40.940 34.620 41.440 34.790 ;
        RECT 41.730 34.620 42.230 34.790 ;
        RECT 42.520 34.620 43.020 34.790 ;
        RECT 45.210 34.620 45.710 34.790 ;
        RECT 46.000 34.620 46.500 34.790 ;
        RECT 46.790 34.620 47.290 34.790 ;
        RECT 47.580 34.620 48.080 34.790 ;
        RECT 48.370 34.620 48.870 34.790 ;
        RECT 49.160 34.620 49.660 34.790 ;
        RECT 49.950 34.620 50.450 34.790 ;
        RECT 50.740 34.620 51.240 34.790 ;
        RECT 51.530 34.620 52.030 34.790 ;
        RECT 52.320 34.620 52.820 34.790 ;
        RECT 55.010 34.620 55.510 34.790 ;
        RECT 55.800 34.620 56.300 34.790 ;
        RECT 56.590 34.620 57.090 34.790 ;
        RECT 57.380 34.620 57.880 34.790 ;
        RECT 58.170 34.620 58.670 34.790 ;
        RECT 58.960 34.620 59.460 34.790 ;
        RECT 59.750 34.620 60.250 34.790 ;
        RECT 60.540 34.620 61.040 34.790 ;
        RECT 61.330 34.620 61.830 34.790 ;
        RECT 62.120 34.620 62.620 34.790 ;
        RECT 64.810 34.620 65.310 34.790 ;
        RECT 65.600 34.620 66.100 34.790 ;
        RECT 66.390 34.620 66.890 34.790 ;
        RECT 67.180 34.620 67.680 34.790 ;
        RECT 67.970 34.620 68.470 34.790 ;
        RECT 68.760 34.620 69.260 34.790 ;
        RECT 69.550 34.620 70.050 34.790 ;
        RECT 70.340 34.620 70.840 34.790 ;
        RECT 71.130 34.620 71.630 34.790 ;
        RECT 71.920 34.620 72.420 34.790 ;
        RECT 25.470 34.080 25.970 34.250 ;
        RECT 26.260 34.080 26.760 34.250 ;
        RECT 27.050 34.080 27.550 34.250 ;
        RECT 27.840 34.080 28.340 34.250 ;
        RECT 28.630 34.080 29.130 34.250 ;
        RECT 29.420 34.080 29.920 34.250 ;
        RECT 30.210 34.080 30.710 34.250 ;
        RECT 31.000 34.080 31.500 34.250 ;
        RECT 31.790 34.080 32.290 34.250 ;
        RECT 32.580 34.080 33.080 34.250 ;
        RECT 35.410 34.080 35.910 34.250 ;
        RECT 36.200 34.080 36.700 34.250 ;
        RECT 36.990 34.080 37.490 34.250 ;
        RECT 37.780 34.080 38.280 34.250 ;
        RECT 38.570 34.080 39.070 34.250 ;
        RECT 39.360 34.080 39.860 34.250 ;
        RECT 40.150 34.080 40.650 34.250 ;
        RECT 40.940 34.080 41.440 34.250 ;
        RECT 41.730 34.080 42.230 34.250 ;
        RECT 42.520 34.080 43.020 34.250 ;
        RECT 45.210 34.080 45.710 34.250 ;
        RECT 46.000 34.080 46.500 34.250 ;
        RECT 46.790 34.080 47.290 34.250 ;
        RECT 47.580 34.080 48.080 34.250 ;
        RECT 48.370 34.080 48.870 34.250 ;
        RECT 49.160 34.080 49.660 34.250 ;
        RECT 49.950 34.080 50.450 34.250 ;
        RECT 50.740 34.080 51.240 34.250 ;
        RECT 51.530 34.080 52.030 34.250 ;
        RECT 52.320 34.080 52.820 34.250 ;
        RECT 55.010 34.080 55.510 34.250 ;
        RECT 55.800 34.080 56.300 34.250 ;
        RECT 56.590 34.080 57.090 34.250 ;
        RECT 57.380 34.080 57.880 34.250 ;
        RECT 58.170 34.080 58.670 34.250 ;
        RECT 58.960 34.080 59.460 34.250 ;
        RECT 59.750 34.080 60.250 34.250 ;
        RECT 60.540 34.080 61.040 34.250 ;
        RECT 61.330 34.080 61.830 34.250 ;
        RECT 62.120 34.080 62.620 34.250 ;
        RECT 64.810 34.080 65.310 34.250 ;
        RECT 65.600 34.080 66.100 34.250 ;
        RECT 66.390 34.080 66.890 34.250 ;
        RECT 67.180 34.080 67.680 34.250 ;
        RECT 67.970 34.080 68.470 34.250 ;
        RECT 68.760 34.080 69.260 34.250 ;
        RECT 69.550 34.080 70.050 34.250 ;
        RECT 70.340 34.080 70.840 34.250 ;
        RECT 71.130 34.080 71.630 34.250 ;
        RECT 71.920 34.080 72.420 34.250 ;
        RECT 16.540 24.840 17.040 25.010 ;
        RECT 17.330 24.840 17.830 25.010 ;
        RECT 20.025 24.835 20.525 25.005 ;
        RECT 20.815 24.835 21.315 25.005 ;
        RECT 21.605 24.835 22.105 25.005 ;
        RECT 22.395 24.835 22.895 25.005 ;
        RECT 25.470 23.440 25.970 23.610 ;
        RECT 26.260 23.440 26.760 23.610 ;
        RECT 27.050 23.440 27.550 23.610 ;
        RECT 27.840 23.440 28.340 23.610 ;
        RECT 28.630 23.440 29.130 23.610 ;
        RECT 29.420 23.440 29.920 23.610 ;
        RECT 30.210 23.440 30.710 23.610 ;
        RECT 31.000 23.440 31.500 23.610 ;
        RECT 31.790 23.440 32.290 23.610 ;
        RECT 32.580 23.440 33.080 23.610 ;
        RECT 35.410 23.440 35.910 23.610 ;
        RECT 36.200 23.440 36.700 23.610 ;
        RECT 36.990 23.440 37.490 23.610 ;
        RECT 37.780 23.440 38.280 23.610 ;
        RECT 38.570 23.440 39.070 23.610 ;
        RECT 39.360 23.440 39.860 23.610 ;
        RECT 40.150 23.440 40.650 23.610 ;
        RECT 40.940 23.440 41.440 23.610 ;
        RECT 41.730 23.440 42.230 23.610 ;
        RECT 42.520 23.440 43.020 23.610 ;
        RECT 45.210 23.440 45.710 23.610 ;
        RECT 46.000 23.440 46.500 23.610 ;
        RECT 46.790 23.440 47.290 23.610 ;
        RECT 47.580 23.440 48.080 23.610 ;
        RECT 48.370 23.440 48.870 23.610 ;
        RECT 49.160 23.440 49.660 23.610 ;
        RECT 49.950 23.440 50.450 23.610 ;
        RECT 50.740 23.440 51.240 23.610 ;
        RECT 51.530 23.440 52.030 23.610 ;
        RECT 52.320 23.440 52.820 23.610 ;
        RECT 55.010 23.440 55.510 23.610 ;
        RECT 55.800 23.440 56.300 23.610 ;
        RECT 56.590 23.440 57.090 23.610 ;
        RECT 57.380 23.440 57.880 23.610 ;
        RECT 58.170 23.440 58.670 23.610 ;
        RECT 58.960 23.440 59.460 23.610 ;
        RECT 59.750 23.440 60.250 23.610 ;
        RECT 60.540 23.440 61.040 23.610 ;
        RECT 61.330 23.440 61.830 23.610 ;
        RECT 62.120 23.440 62.620 23.610 ;
        RECT 64.810 23.440 65.310 23.610 ;
        RECT 65.600 23.440 66.100 23.610 ;
        RECT 66.390 23.440 66.890 23.610 ;
        RECT 67.180 23.440 67.680 23.610 ;
        RECT 67.970 23.440 68.470 23.610 ;
        RECT 68.760 23.440 69.260 23.610 ;
        RECT 69.550 23.440 70.050 23.610 ;
        RECT 70.340 23.440 70.840 23.610 ;
        RECT 71.130 23.440 71.630 23.610 ;
        RECT 71.920 23.440 72.420 23.610 ;
        RECT 15.285 22.905 15.785 23.075 ;
        RECT 16.075 22.905 16.575 23.075 ;
        RECT 16.865 22.905 17.365 23.075 ;
        RECT 17.655 22.905 18.155 23.075 ;
        RECT 18.445 22.905 18.945 23.075 ;
        RECT 19.235 22.905 19.735 23.075 ;
        RECT 20.025 22.905 20.525 23.075 ;
        RECT 20.815 22.905 21.315 23.075 ;
        RECT 21.605 22.905 22.105 23.075 ;
        RECT 22.395 22.905 22.895 23.075 ;
        RECT 25.470 22.900 25.970 23.070 ;
        RECT 26.260 22.900 26.760 23.070 ;
        RECT 27.050 22.900 27.550 23.070 ;
        RECT 27.840 22.900 28.340 23.070 ;
        RECT 28.630 22.900 29.130 23.070 ;
        RECT 29.420 22.900 29.920 23.070 ;
        RECT 30.210 22.900 30.710 23.070 ;
        RECT 31.000 22.900 31.500 23.070 ;
        RECT 31.790 22.900 32.290 23.070 ;
        RECT 32.580 22.900 33.080 23.070 ;
        RECT 35.410 22.900 35.910 23.070 ;
        RECT 36.200 22.900 36.700 23.070 ;
        RECT 36.990 22.900 37.490 23.070 ;
        RECT 37.780 22.900 38.280 23.070 ;
        RECT 38.570 22.900 39.070 23.070 ;
        RECT 39.360 22.900 39.860 23.070 ;
        RECT 40.150 22.900 40.650 23.070 ;
        RECT 40.940 22.900 41.440 23.070 ;
        RECT 41.730 22.900 42.230 23.070 ;
        RECT 42.520 22.900 43.020 23.070 ;
        RECT 45.210 22.900 45.710 23.070 ;
        RECT 46.000 22.900 46.500 23.070 ;
        RECT 46.790 22.900 47.290 23.070 ;
        RECT 47.580 22.900 48.080 23.070 ;
        RECT 48.370 22.900 48.870 23.070 ;
        RECT 49.160 22.900 49.660 23.070 ;
        RECT 49.950 22.900 50.450 23.070 ;
        RECT 50.740 22.900 51.240 23.070 ;
        RECT 51.530 22.900 52.030 23.070 ;
        RECT 52.320 22.900 52.820 23.070 ;
        RECT 55.010 22.900 55.510 23.070 ;
        RECT 55.800 22.900 56.300 23.070 ;
        RECT 56.590 22.900 57.090 23.070 ;
        RECT 57.380 22.900 57.880 23.070 ;
        RECT 58.170 22.900 58.670 23.070 ;
        RECT 58.960 22.900 59.460 23.070 ;
        RECT 59.750 22.900 60.250 23.070 ;
        RECT 60.540 22.900 61.040 23.070 ;
        RECT 61.330 22.900 61.830 23.070 ;
        RECT 62.120 22.900 62.620 23.070 ;
        RECT 64.810 22.900 65.310 23.070 ;
        RECT 65.600 22.900 66.100 23.070 ;
        RECT 66.390 22.900 66.890 23.070 ;
        RECT 67.180 22.900 67.680 23.070 ;
        RECT 67.970 22.900 68.470 23.070 ;
        RECT 68.760 22.900 69.260 23.070 ;
        RECT 69.550 22.900 70.050 23.070 ;
        RECT 70.340 22.900 70.840 23.070 ;
        RECT 71.130 22.900 71.630 23.070 ;
        RECT 71.920 22.900 72.420 23.070 ;
        RECT 15.845 12.645 16.015 22.685 ;
        RECT 17.425 12.645 17.595 22.685 ;
        RECT 19.005 12.645 19.175 22.685 ;
        RECT 20.585 12.645 20.755 22.685 ;
        RECT 22.165 12.645 22.335 22.685 ;
        RECT 15.285 12.255 15.785 12.425 ;
        RECT 16.075 12.255 16.575 12.425 ;
        RECT 16.865 12.255 17.365 12.425 ;
        RECT 17.655 12.255 18.155 12.425 ;
        RECT 18.445 12.255 18.945 12.425 ;
        RECT 19.235 12.255 19.735 12.425 ;
        RECT 20.025 12.255 20.525 12.425 ;
        RECT 20.815 12.255 21.315 12.425 ;
        RECT 21.605 12.255 22.105 12.425 ;
        RECT 22.395 12.255 22.895 12.425 ;
        RECT 25.470 12.260 25.970 12.430 ;
        RECT 26.260 12.260 26.760 12.430 ;
        RECT 27.050 12.260 27.550 12.430 ;
        RECT 27.840 12.260 28.340 12.430 ;
        RECT 28.630 12.260 29.130 12.430 ;
        RECT 29.420 12.260 29.920 12.430 ;
        RECT 30.210 12.260 30.710 12.430 ;
        RECT 31.000 12.260 31.500 12.430 ;
        RECT 31.790 12.260 32.290 12.430 ;
        RECT 32.580 12.260 33.080 12.430 ;
        RECT 35.410 12.260 35.910 12.430 ;
        RECT 36.200 12.260 36.700 12.430 ;
        RECT 36.990 12.260 37.490 12.430 ;
        RECT 37.780 12.260 38.280 12.430 ;
        RECT 38.570 12.260 39.070 12.430 ;
        RECT 39.360 12.260 39.860 12.430 ;
        RECT 40.150 12.260 40.650 12.430 ;
        RECT 40.940 12.260 41.440 12.430 ;
        RECT 41.730 12.260 42.230 12.430 ;
        RECT 42.520 12.260 43.020 12.430 ;
        RECT 45.210 12.260 45.710 12.430 ;
        RECT 46.000 12.260 46.500 12.430 ;
        RECT 46.790 12.260 47.290 12.430 ;
        RECT 47.580 12.260 48.080 12.430 ;
        RECT 48.370 12.260 48.870 12.430 ;
        RECT 49.160 12.260 49.660 12.430 ;
        RECT 49.950 12.260 50.450 12.430 ;
        RECT 50.740 12.260 51.240 12.430 ;
        RECT 51.530 12.260 52.030 12.430 ;
        RECT 52.320 12.260 52.820 12.430 ;
        RECT 55.010 12.260 55.510 12.430 ;
        RECT 55.800 12.260 56.300 12.430 ;
        RECT 56.590 12.260 57.090 12.430 ;
        RECT 57.380 12.260 57.880 12.430 ;
        RECT 58.170 12.260 58.670 12.430 ;
        RECT 58.960 12.260 59.460 12.430 ;
        RECT 59.750 12.260 60.250 12.430 ;
        RECT 60.540 12.260 61.040 12.430 ;
        RECT 61.330 12.260 61.830 12.430 ;
        RECT 62.120 12.260 62.620 12.430 ;
        RECT 64.810 12.260 65.310 12.430 ;
        RECT 65.600 12.260 66.100 12.430 ;
        RECT 66.390 12.260 66.890 12.430 ;
        RECT 67.180 12.260 67.680 12.430 ;
        RECT 67.970 12.260 68.470 12.430 ;
        RECT 68.760 12.260 69.260 12.430 ;
        RECT 69.550 12.260 70.050 12.430 ;
        RECT 70.340 12.260 70.840 12.430 ;
        RECT 71.130 12.260 71.630 12.430 ;
        RECT 71.920 12.260 72.420 12.430 ;
        RECT 15.285 11.725 15.785 11.895 ;
        RECT 16.075 11.725 16.575 11.895 ;
        RECT 16.865 11.725 17.365 11.895 ;
        RECT 17.655 11.725 18.155 11.895 ;
        RECT 18.445 11.725 18.945 11.895 ;
        RECT 19.235 11.725 19.735 11.895 ;
        RECT 20.025 11.725 20.525 11.895 ;
        RECT 20.815 11.725 21.315 11.895 ;
        RECT 21.605 11.725 22.105 11.895 ;
        RECT 22.395 11.725 22.895 11.895 ;
        RECT 25.470 11.720 25.970 11.890 ;
        RECT 26.260 11.720 26.760 11.890 ;
        RECT 27.050 11.720 27.550 11.890 ;
        RECT 27.840 11.720 28.340 11.890 ;
        RECT 28.630 11.720 29.130 11.890 ;
        RECT 29.420 11.720 29.920 11.890 ;
        RECT 30.210 11.720 30.710 11.890 ;
        RECT 31.000 11.720 31.500 11.890 ;
        RECT 31.790 11.720 32.290 11.890 ;
        RECT 32.580 11.720 33.080 11.890 ;
        RECT 35.410 11.720 35.910 11.890 ;
        RECT 36.200 11.720 36.700 11.890 ;
        RECT 36.990 11.720 37.490 11.890 ;
        RECT 37.780 11.720 38.280 11.890 ;
        RECT 38.570 11.720 39.070 11.890 ;
        RECT 39.360 11.720 39.860 11.890 ;
        RECT 40.150 11.720 40.650 11.890 ;
        RECT 40.940 11.720 41.440 11.890 ;
        RECT 41.730 11.720 42.230 11.890 ;
        RECT 42.520 11.720 43.020 11.890 ;
        RECT 45.210 11.720 45.710 11.890 ;
        RECT 46.000 11.720 46.500 11.890 ;
        RECT 46.790 11.720 47.290 11.890 ;
        RECT 47.580 11.720 48.080 11.890 ;
        RECT 48.370 11.720 48.870 11.890 ;
        RECT 49.160 11.720 49.660 11.890 ;
        RECT 49.950 11.720 50.450 11.890 ;
        RECT 50.740 11.720 51.240 11.890 ;
        RECT 51.530 11.720 52.030 11.890 ;
        RECT 52.320 11.720 52.820 11.890 ;
        RECT 55.010 11.720 55.510 11.890 ;
        RECT 55.800 11.720 56.300 11.890 ;
        RECT 56.590 11.720 57.090 11.890 ;
        RECT 57.380 11.720 57.880 11.890 ;
        RECT 58.170 11.720 58.670 11.890 ;
        RECT 58.960 11.720 59.460 11.890 ;
        RECT 59.750 11.720 60.250 11.890 ;
        RECT 60.540 11.720 61.040 11.890 ;
        RECT 61.330 11.720 61.830 11.890 ;
        RECT 62.120 11.720 62.620 11.890 ;
        RECT 64.810 11.720 65.310 11.890 ;
        RECT 65.600 11.720 66.100 11.890 ;
        RECT 66.390 11.720 66.890 11.890 ;
        RECT 67.180 11.720 67.680 11.890 ;
        RECT 67.970 11.720 68.470 11.890 ;
        RECT 68.760 11.720 69.260 11.890 ;
        RECT 69.550 11.720 70.050 11.890 ;
        RECT 70.340 11.720 70.840 11.890 ;
        RECT 71.130 11.720 71.630 11.890 ;
        RECT 71.920 11.720 72.420 11.890 ;
        RECT 15.845 1.465 16.015 11.505 ;
        RECT 17.425 1.465 17.595 11.505 ;
        RECT 19.005 1.465 19.175 11.505 ;
        RECT 20.585 1.465 20.755 11.505 ;
        RECT 22.165 1.465 22.335 11.505 ;
        RECT 15.285 1.075 15.785 1.245 ;
        RECT 16.075 1.075 16.575 1.245 ;
        RECT 16.865 1.075 17.365 1.245 ;
        RECT 17.655 1.075 18.155 1.245 ;
        RECT 18.445 1.075 18.945 1.245 ;
        RECT 19.235 1.075 19.735 1.245 ;
        RECT 20.025 1.075 20.525 1.245 ;
        RECT 20.815 1.075 21.315 1.245 ;
        RECT 21.605 1.075 22.105 1.245 ;
        RECT 22.395 1.075 22.895 1.245 ;
        RECT 25.470 1.080 25.970 1.250 ;
        RECT 26.260 1.080 26.760 1.250 ;
        RECT 27.050 1.080 27.550 1.250 ;
        RECT 27.840 1.080 28.340 1.250 ;
        RECT 28.630 1.080 29.130 1.250 ;
        RECT 29.420 1.080 29.920 1.250 ;
        RECT 30.210 1.080 30.710 1.250 ;
        RECT 31.000 1.080 31.500 1.250 ;
        RECT 31.790 1.080 32.290 1.250 ;
        RECT 32.580 1.080 33.080 1.250 ;
        RECT 35.410 1.080 35.910 1.250 ;
        RECT 36.200 1.080 36.700 1.250 ;
        RECT 36.990 1.080 37.490 1.250 ;
        RECT 37.780 1.080 38.280 1.250 ;
        RECT 38.570 1.080 39.070 1.250 ;
        RECT 39.360 1.080 39.860 1.250 ;
        RECT 40.150 1.080 40.650 1.250 ;
        RECT 40.940 1.080 41.440 1.250 ;
        RECT 41.730 1.080 42.230 1.250 ;
        RECT 42.520 1.080 43.020 1.250 ;
        RECT 45.210 1.080 45.710 1.250 ;
        RECT 46.000 1.080 46.500 1.250 ;
        RECT 46.790 1.080 47.290 1.250 ;
        RECT 47.580 1.080 48.080 1.250 ;
        RECT 48.370 1.080 48.870 1.250 ;
        RECT 49.160 1.080 49.660 1.250 ;
        RECT 49.950 1.080 50.450 1.250 ;
        RECT 50.740 1.080 51.240 1.250 ;
        RECT 51.530 1.080 52.030 1.250 ;
        RECT 52.320 1.080 52.820 1.250 ;
        RECT 55.010 1.080 55.510 1.250 ;
        RECT 55.800 1.080 56.300 1.250 ;
        RECT 56.590 1.080 57.090 1.250 ;
        RECT 57.380 1.080 57.880 1.250 ;
        RECT 58.170 1.080 58.670 1.250 ;
        RECT 58.960 1.080 59.460 1.250 ;
        RECT 59.750 1.080 60.250 1.250 ;
        RECT 60.540 1.080 61.040 1.250 ;
        RECT 61.330 1.080 61.830 1.250 ;
        RECT 62.120 1.080 62.620 1.250 ;
        RECT 64.810 1.080 65.310 1.250 ;
        RECT 65.600 1.080 66.100 1.250 ;
        RECT 66.390 1.080 66.890 1.250 ;
        RECT 67.180 1.080 67.680 1.250 ;
        RECT 67.970 1.080 68.470 1.250 ;
        RECT 68.760 1.080 69.260 1.250 ;
        RECT 69.550 1.080 70.050 1.250 ;
        RECT 70.340 1.080 70.840 1.250 ;
        RECT 71.130 1.080 71.630 1.250 ;
        RECT 71.920 1.080 72.420 1.250 ;
      LAYER mcon ;
        RECT 15.365 140.585 15.705 140.755 ;
        RECT 16.155 140.585 16.495 140.755 ;
        RECT 16.945 140.585 17.285 140.755 ;
        RECT 17.735 140.585 18.075 140.755 ;
        RECT 18.525 140.585 18.865 140.755 ;
        RECT 19.315 140.585 19.655 140.755 ;
        RECT 20.105 140.585 20.445 140.755 ;
        RECT 20.895 140.585 21.235 140.755 ;
        RECT 21.685 140.585 22.025 140.755 ;
        RECT 22.475 140.585 22.815 140.755 ;
        RECT 25.550 140.580 25.890 140.750 ;
        RECT 26.340 140.580 26.680 140.750 ;
        RECT 27.130 140.580 27.470 140.750 ;
        RECT 27.920 140.580 28.260 140.750 ;
        RECT 28.710 140.580 29.050 140.750 ;
        RECT 29.500 140.580 29.840 140.750 ;
        RECT 30.290 140.580 30.630 140.750 ;
        RECT 31.080 140.580 31.420 140.750 ;
        RECT 31.870 140.580 32.210 140.750 ;
        RECT 32.660 140.580 33.000 140.750 ;
        RECT 35.490 140.580 35.830 140.750 ;
        RECT 36.280 140.580 36.620 140.750 ;
        RECT 37.070 140.580 37.410 140.750 ;
        RECT 37.860 140.580 38.200 140.750 ;
        RECT 38.650 140.580 38.990 140.750 ;
        RECT 39.440 140.580 39.780 140.750 ;
        RECT 40.230 140.580 40.570 140.750 ;
        RECT 41.020 140.580 41.360 140.750 ;
        RECT 41.810 140.580 42.150 140.750 ;
        RECT 42.600 140.580 42.940 140.750 ;
        RECT 45.290 140.580 45.630 140.750 ;
        RECT 46.080 140.580 46.420 140.750 ;
        RECT 46.870 140.580 47.210 140.750 ;
        RECT 47.660 140.580 48.000 140.750 ;
        RECT 48.450 140.580 48.790 140.750 ;
        RECT 49.240 140.580 49.580 140.750 ;
        RECT 50.030 140.580 50.370 140.750 ;
        RECT 50.820 140.580 51.160 140.750 ;
        RECT 51.610 140.580 51.950 140.750 ;
        RECT 52.400 140.580 52.740 140.750 ;
        RECT 55.090 140.580 55.430 140.750 ;
        RECT 55.880 140.580 56.220 140.750 ;
        RECT 56.670 140.580 57.010 140.750 ;
        RECT 57.460 140.580 57.800 140.750 ;
        RECT 58.250 140.580 58.590 140.750 ;
        RECT 59.040 140.580 59.380 140.750 ;
        RECT 59.830 140.580 60.170 140.750 ;
        RECT 60.620 140.580 60.960 140.750 ;
        RECT 61.410 140.580 61.750 140.750 ;
        RECT 62.200 140.580 62.540 140.750 ;
        RECT 64.890 140.580 65.230 140.750 ;
        RECT 65.680 140.580 66.020 140.750 ;
        RECT 66.470 140.580 66.810 140.750 ;
        RECT 67.260 140.580 67.600 140.750 ;
        RECT 68.050 140.580 68.390 140.750 ;
        RECT 68.840 140.580 69.180 140.750 ;
        RECT 69.630 140.580 69.970 140.750 ;
        RECT 70.420 140.580 70.760 140.750 ;
        RECT 71.210 140.580 71.550 140.750 ;
        RECT 72.000 140.580 72.340 140.750 ;
        RECT 15.845 130.405 16.015 140.285 ;
        RECT 17.425 130.405 17.595 140.285 ;
        RECT 19.005 130.405 19.175 140.285 ;
        RECT 20.585 130.405 20.755 140.285 ;
        RECT 22.165 130.405 22.335 140.285 ;
        RECT 15.365 129.935 15.705 130.105 ;
        RECT 16.155 129.935 16.495 130.105 ;
        RECT 16.945 129.935 17.285 130.105 ;
        RECT 17.735 129.935 18.075 130.105 ;
        RECT 18.525 129.935 18.865 130.105 ;
        RECT 19.315 129.935 19.655 130.105 ;
        RECT 20.105 129.935 20.445 130.105 ;
        RECT 20.895 129.935 21.235 130.105 ;
        RECT 21.685 129.935 22.025 130.105 ;
        RECT 22.475 129.935 22.815 130.105 ;
        RECT 25.550 129.940 25.890 130.110 ;
        RECT 26.340 129.940 26.680 130.110 ;
        RECT 27.130 129.940 27.470 130.110 ;
        RECT 27.920 129.940 28.260 130.110 ;
        RECT 28.710 129.940 29.050 130.110 ;
        RECT 29.500 129.940 29.840 130.110 ;
        RECT 30.290 129.940 30.630 130.110 ;
        RECT 31.080 129.940 31.420 130.110 ;
        RECT 31.870 129.940 32.210 130.110 ;
        RECT 32.660 129.940 33.000 130.110 ;
        RECT 35.490 129.940 35.830 130.110 ;
        RECT 36.280 129.940 36.620 130.110 ;
        RECT 37.070 129.940 37.410 130.110 ;
        RECT 37.860 129.940 38.200 130.110 ;
        RECT 38.650 129.940 38.990 130.110 ;
        RECT 39.440 129.940 39.780 130.110 ;
        RECT 40.230 129.940 40.570 130.110 ;
        RECT 41.020 129.940 41.360 130.110 ;
        RECT 41.810 129.940 42.150 130.110 ;
        RECT 42.600 129.940 42.940 130.110 ;
        RECT 45.290 129.940 45.630 130.110 ;
        RECT 46.080 129.940 46.420 130.110 ;
        RECT 46.870 129.940 47.210 130.110 ;
        RECT 47.660 129.940 48.000 130.110 ;
        RECT 48.450 129.940 48.790 130.110 ;
        RECT 49.240 129.940 49.580 130.110 ;
        RECT 50.030 129.940 50.370 130.110 ;
        RECT 50.820 129.940 51.160 130.110 ;
        RECT 51.610 129.940 51.950 130.110 ;
        RECT 52.400 129.940 52.740 130.110 ;
        RECT 55.090 129.940 55.430 130.110 ;
        RECT 55.880 129.940 56.220 130.110 ;
        RECT 56.670 129.940 57.010 130.110 ;
        RECT 57.460 129.940 57.800 130.110 ;
        RECT 58.250 129.940 58.590 130.110 ;
        RECT 59.040 129.940 59.380 130.110 ;
        RECT 59.830 129.940 60.170 130.110 ;
        RECT 60.620 129.940 60.960 130.110 ;
        RECT 61.410 129.940 61.750 130.110 ;
        RECT 62.200 129.940 62.540 130.110 ;
        RECT 64.890 129.940 65.230 130.110 ;
        RECT 65.680 129.940 66.020 130.110 ;
        RECT 66.470 129.940 66.810 130.110 ;
        RECT 67.260 129.940 67.600 130.110 ;
        RECT 68.050 129.940 68.390 130.110 ;
        RECT 68.840 129.940 69.180 130.110 ;
        RECT 69.630 129.940 69.970 130.110 ;
        RECT 70.420 129.940 70.760 130.110 ;
        RECT 71.210 129.940 71.550 130.110 ;
        RECT 72.000 129.940 72.340 130.110 ;
        RECT 15.365 129.405 15.705 129.575 ;
        RECT 16.155 129.405 16.495 129.575 ;
        RECT 16.945 129.405 17.285 129.575 ;
        RECT 17.735 129.405 18.075 129.575 ;
        RECT 18.525 129.405 18.865 129.575 ;
        RECT 19.315 129.405 19.655 129.575 ;
        RECT 20.105 129.405 20.445 129.575 ;
        RECT 20.895 129.405 21.235 129.575 ;
        RECT 21.685 129.405 22.025 129.575 ;
        RECT 22.475 129.405 22.815 129.575 ;
        RECT 25.550 129.400 25.890 129.570 ;
        RECT 26.340 129.400 26.680 129.570 ;
        RECT 27.130 129.400 27.470 129.570 ;
        RECT 27.920 129.400 28.260 129.570 ;
        RECT 28.710 129.400 29.050 129.570 ;
        RECT 29.500 129.400 29.840 129.570 ;
        RECT 30.290 129.400 30.630 129.570 ;
        RECT 31.080 129.400 31.420 129.570 ;
        RECT 31.870 129.400 32.210 129.570 ;
        RECT 32.660 129.400 33.000 129.570 ;
        RECT 35.490 129.400 35.830 129.570 ;
        RECT 36.280 129.400 36.620 129.570 ;
        RECT 37.070 129.400 37.410 129.570 ;
        RECT 37.860 129.400 38.200 129.570 ;
        RECT 38.650 129.400 38.990 129.570 ;
        RECT 39.440 129.400 39.780 129.570 ;
        RECT 40.230 129.400 40.570 129.570 ;
        RECT 41.020 129.400 41.360 129.570 ;
        RECT 41.810 129.400 42.150 129.570 ;
        RECT 42.600 129.400 42.940 129.570 ;
        RECT 45.290 129.400 45.630 129.570 ;
        RECT 46.080 129.400 46.420 129.570 ;
        RECT 46.870 129.400 47.210 129.570 ;
        RECT 47.660 129.400 48.000 129.570 ;
        RECT 48.450 129.400 48.790 129.570 ;
        RECT 49.240 129.400 49.580 129.570 ;
        RECT 50.030 129.400 50.370 129.570 ;
        RECT 50.820 129.400 51.160 129.570 ;
        RECT 51.610 129.400 51.950 129.570 ;
        RECT 52.400 129.400 52.740 129.570 ;
        RECT 55.090 129.400 55.430 129.570 ;
        RECT 55.880 129.400 56.220 129.570 ;
        RECT 56.670 129.400 57.010 129.570 ;
        RECT 57.460 129.400 57.800 129.570 ;
        RECT 58.250 129.400 58.590 129.570 ;
        RECT 59.040 129.400 59.380 129.570 ;
        RECT 59.830 129.400 60.170 129.570 ;
        RECT 60.620 129.400 60.960 129.570 ;
        RECT 61.410 129.400 61.750 129.570 ;
        RECT 62.200 129.400 62.540 129.570 ;
        RECT 64.890 129.400 65.230 129.570 ;
        RECT 65.680 129.400 66.020 129.570 ;
        RECT 66.470 129.400 66.810 129.570 ;
        RECT 67.260 129.400 67.600 129.570 ;
        RECT 68.050 129.400 68.390 129.570 ;
        RECT 68.840 129.400 69.180 129.570 ;
        RECT 69.630 129.400 69.970 129.570 ;
        RECT 70.420 129.400 70.760 129.570 ;
        RECT 71.210 129.400 71.550 129.570 ;
        RECT 72.000 129.400 72.340 129.570 ;
        RECT 15.845 119.225 16.015 129.105 ;
        RECT 17.425 119.225 17.595 129.105 ;
        RECT 19.005 119.225 19.175 129.105 ;
        RECT 20.585 119.225 20.755 129.105 ;
        RECT 22.165 119.225 22.335 129.105 ;
        RECT 15.365 118.755 15.705 118.925 ;
        RECT 16.155 118.755 16.495 118.925 ;
        RECT 16.945 118.755 17.285 118.925 ;
        RECT 17.735 118.755 18.075 118.925 ;
        RECT 18.525 118.755 18.865 118.925 ;
        RECT 19.315 118.755 19.655 118.925 ;
        RECT 20.105 118.755 20.445 118.925 ;
        RECT 20.895 118.755 21.235 118.925 ;
        RECT 21.685 118.755 22.025 118.925 ;
        RECT 22.475 118.755 22.815 118.925 ;
        RECT 25.550 118.760 25.890 118.930 ;
        RECT 26.340 118.760 26.680 118.930 ;
        RECT 27.130 118.760 27.470 118.930 ;
        RECT 27.920 118.760 28.260 118.930 ;
        RECT 28.710 118.760 29.050 118.930 ;
        RECT 29.500 118.760 29.840 118.930 ;
        RECT 30.290 118.760 30.630 118.930 ;
        RECT 31.080 118.760 31.420 118.930 ;
        RECT 31.870 118.760 32.210 118.930 ;
        RECT 32.660 118.760 33.000 118.930 ;
        RECT 35.490 118.760 35.830 118.930 ;
        RECT 36.280 118.760 36.620 118.930 ;
        RECT 37.070 118.760 37.410 118.930 ;
        RECT 37.860 118.760 38.200 118.930 ;
        RECT 38.650 118.760 38.990 118.930 ;
        RECT 39.440 118.760 39.780 118.930 ;
        RECT 40.230 118.760 40.570 118.930 ;
        RECT 41.020 118.760 41.360 118.930 ;
        RECT 41.810 118.760 42.150 118.930 ;
        RECT 42.600 118.760 42.940 118.930 ;
        RECT 45.290 118.760 45.630 118.930 ;
        RECT 46.080 118.760 46.420 118.930 ;
        RECT 46.870 118.760 47.210 118.930 ;
        RECT 47.660 118.760 48.000 118.930 ;
        RECT 48.450 118.760 48.790 118.930 ;
        RECT 49.240 118.760 49.580 118.930 ;
        RECT 50.030 118.760 50.370 118.930 ;
        RECT 50.820 118.760 51.160 118.930 ;
        RECT 51.610 118.760 51.950 118.930 ;
        RECT 52.400 118.760 52.740 118.930 ;
        RECT 55.090 118.760 55.430 118.930 ;
        RECT 55.880 118.760 56.220 118.930 ;
        RECT 56.670 118.760 57.010 118.930 ;
        RECT 57.460 118.760 57.800 118.930 ;
        RECT 58.250 118.760 58.590 118.930 ;
        RECT 59.040 118.760 59.380 118.930 ;
        RECT 59.830 118.760 60.170 118.930 ;
        RECT 60.620 118.760 60.960 118.930 ;
        RECT 61.410 118.760 61.750 118.930 ;
        RECT 62.200 118.760 62.540 118.930 ;
        RECT 64.890 118.760 65.230 118.930 ;
        RECT 65.680 118.760 66.020 118.930 ;
        RECT 66.470 118.760 66.810 118.930 ;
        RECT 67.260 118.760 67.600 118.930 ;
        RECT 68.050 118.760 68.390 118.930 ;
        RECT 68.840 118.760 69.180 118.930 ;
        RECT 69.630 118.760 69.970 118.930 ;
        RECT 70.420 118.760 70.760 118.930 ;
        RECT 71.210 118.760 71.550 118.930 ;
        RECT 72.000 118.760 72.340 118.930 ;
        RECT 25.550 118.220 25.890 118.390 ;
        RECT 26.340 118.220 26.680 118.390 ;
        RECT 27.130 118.220 27.470 118.390 ;
        RECT 27.920 118.220 28.260 118.390 ;
        RECT 28.710 118.220 29.050 118.390 ;
        RECT 29.500 118.220 29.840 118.390 ;
        RECT 30.290 118.220 30.630 118.390 ;
        RECT 31.080 118.220 31.420 118.390 ;
        RECT 31.870 118.220 32.210 118.390 ;
        RECT 32.660 118.220 33.000 118.390 ;
        RECT 35.490 118.220 35.830 118.390 ;
        RECT 36.280 118.220 36.620 118.390 ;
        RECT 37.070 118.220 37.410 118.390 ;
        RECT 37.860 118.220 38.200 118.390 ;
        RECT 38.650 118.220 38.990 118.390 ;
        RECT 39.440 118.220 39.780 118.390 ;
        RECT 40.230 118.220 40.570 118.390 ;
        RECT 41.020 118.220 41.360 118.390 ;
        RECT 41.810 118.220 42.150 118.390 ;
        RECT 42.600 118.220 42.940 118.390 ;
        RECT 45.290 118.220 45.630 118.390 ;
        RECT 46.080 118.220 46.420 118.390 ;
        RECT 46.870 118.220 47.210 118.390 ;
        RECT 47.660 118.220 48.000 118.390 ;
        RECT 48.450 118.220 48.790 118.390 ;
        RECT 49.240 118.220 49.580 118.390 ;
        RECT 50.030 118.220 50.370 118.390 ;
        RECT 50.820 118.220 51.160 118.390 ;
        RECT 51.610 118.220 51.950 118.390 ;
        RECT 52.400 118.220 52.740 118.390 ;
        RECT 55.090 118.220 55.430 118.390 ;
        RECT 55.880 118.220 56.220 118.390 ;
        RECT 56.670 118.220 57.010 118.390 ;
        RECT 57.460 118.220 57.800 118.390 ;
        RECT 58.250 118.220 58.590 118.390 ;
        RECT 59.040 118.220 59.380 118.390 ;
        RECT 59.830 118.220 60.170 118.390 ;
        RECT 60.620 118.220 60.960 118.390 ;
        RECT 61.410 118.220 61.750 118.390 ;
        RECT 62.200 118.220 62.540 118.390 ;
        RECT 64.890 118.220 65.230 118.390 ;
        RECT 65.680 118.220 66.020 118.390 ;
        RECT 66.470 118.220 66.810 118.390 ;
        RECT 67.260 118.220 67.600 118.390 ;
        RECT 68.050 118.220 68.390 118.390 ;
        RECT 68.840 118.220 69.180 118.390 ;
        RECT 69.630 118.220 69.970 118.390 ;
        RECT 70.420 118.220 70.760 118.390 ;
        RECT 71.210 118.220 71.550 118.390 ;
        RECT 72.000 118.220 72.340 118.390 ;
        RECT 16.620 116.820 16.960 116.990 ;
        RECT 17.410 116.820 17.750 116.990 ;
        RECT 20.105 116.825 20.445 116.995 ;
        RECT 20.895 116.825 21.235 116.995 ;
        RECT 21.685 116.825 22.025 116.995 ;
        RECT 22.475 116.825 22.815 116.995 ;
        RECT 17.100 112.640 17.270 116.520 ;
        RECT 16.620 112.170 16.960 112.340 ;
        RECT 17.410 112.170 17.750 112.340 ;
        RECT 16.305 109.080 16.475 109.960 ;
        RECT 17.885 109.080 18.055 109.960 ;
        RECT 16.615 108.610 16.955 108.780 ;
        RECT 17.405 108.610 17.745 108.780 ;
        RECT 20.585 106.645 20.755 116.525 ;
        RECT 22.165 106.645 22.335 116.525 ;
        RECT 25.550 107.580 25.890 107.750 ;
        RECT 26.340 107.580 26.680 107.750 ;
        RECT 27.130 107.580 27.470 107.750 ;
        RECT 27.920 107.580 28.260 107.750 ;
        RECT 28.710 107.580 29.050 107.750 ;
        RECT 29.500 107.580 29.840 107.750 ;
        RECT 30.290 107.580 30.630 107.750 ;
        RECT 31.080 107.580 31.420 107.750 ;
        RECT 31.870 107.580 32.210 107.750 ;
        RECT 32.660 107.580 33.000 107.750 ;
        RECT 35.490 107.580 35.830 107.750 ;
        RECT 36.280 107.580 36.620 107.750 ;
        RECT 37.070 107.580 37.410 107.750 ;
        RECT 37.860 107.580 38.200 107.750 ;
        RECT 38.650 107.580 38.990 107.750 ;
        RECT 39.440 107.580 39.780 107.750 ;
        RECT 40.230 107.580 40.570 107.750 ;
        RECT 41.020 107.580 41.360 107.750 ;
        RECT 41.810 107.580 42.150 107.750 ;
        RECT 42.600 107.580 42.940 107.750 ;
        RECT 45.290 107.580 45.630 107.750 ;
        RECT 46.080 107.580 46.420 107.750 ;
        RECT 46.870 107.580 47.210 107.750 ;
        RECT 47.660 107.580 48.000 107.750 ;
        RECT 48.450 107.580 48.790 107.750 ;
        RECT 49.240 107.580 49.580 107.750 ;
        RECT 50.030 107.580 50.370 107.750 ;
        RECT 50.820 107.580 51.160 107.750 ;
        RECT 51.610 107.580 51.950 107.750 ;
        RECT 52.400 107.580 52.740 107.750 ;
        RECT 55.090 107.580 55.430 107.750 ;
        RECT 55.880 107.580 56.220 107.750 ;
        RECT 56.670 107.580 57.010 107.750 ;
        RECT 57.460 107.580 57.800 107.750 ;
        RECT 58.250 107.580 58.590 107.750 ;
        RECT 59.040 107.580 59.380 107.750 ;
        RECT 59.830 107.580 60.170 107.750 ;
        RECT 60.620 107.580 60.960 107.750 ;
        RECT 61.410 107.580 61.750 107.750 ;
        RECT 62.200 107.580 62.540 107.750 ;
        RECT 64.890 107.580 65.230 107.750 ;
        RECT 65.680 107.580 66.020 107.750 ;
        RECT 66.470 107.580 66.810 107.750 ;
        RECT 67.260 107.580 67.600 107.750 ;
        RECT 68.050 107.580 68.390 107.750 ;
        RECT 68.840 107.580 69.180 107.750 ;
        RECT 69.630 107.580 69.970 107.750 ;
        RECT 70.420 107.580 70.760 107.750 ;
        RECT 71.210 107.580 71.550 107.750 ;
        RECT 72.000 107.580 72.340 107.750 ;
        RECT 25.550 107.040 25.890 107.210 ;
        RECT 26.340 107.040 26.680 107.210 ;
        RECT 27.130 107.040 27.470 107.210 ;
        RECT 27.920 107.040 28.260 107.210 ;
        RECT 28.710 107.040 29.050 107.210 ;
        RECT 29.500 107.040 29.840 107.210 ;
        RECT 30.290 107.040 30.630 107.210 ;
        RECT 31.080 107.040 31.420 107.210 ;
        RECT 31.870 107.040 32.210 107.210 ;
        RECT 32.660 107.040 33.000 107.210 ;
        RECT 35.490 107.040 35.830 107.210 ;
        RECT 36.280 107.040 36.620 107.210 ;
        RECT 37.070 107.040 37.410 107.210 ;
        RECT 37.860 107.040 38.200 107.210 ;
        RECT 38.650 107.040 38.990 107.210 ;
        RECT 39.440 107.040 39.780 107.210 ;
        RECT 40.230 107.040 40.570 107.210 ;
        RECT 41.020 107.040 41.360 107.210 ;
        RECT 41.810 107.040 42.150 107.210 ;
        RECT 42.600 107.040 42.940 107.210 ;
        RECT 45.290 107.040 45.630 107.210 ;
        RECT 46.080 107.040 46.420 107.210 ;
        RECT 46.870 107.040 47.210 107.210 ;
        RECT 47.660 107.040 48.000 107.210 ;
        RECT 48.450 107.040 48.790 107.210 ;
        RECT 49.240 107.040 49.580 107.210 ;
        RECT 50.030 107.040 50.370 107.210 ;
        RECT 50.820 107.040 51.160 107.210 ;
        RECT 51.610 107.040 51.950 107.210 ;
        RECT 52.400 107.040 52.740 107.210 ;
        RECT 55.090 107.040 55.430 107.210 ;
        RECT 55.880 107.040 56.220 107.210 ;
        RECT 56.670 107.040 57.010 107.210 ;
        RECT 57.460 107.040 57.800 107.210 ;
        RECT 58.250 107.040 58.590 107.210 ;
        RECT 59.040 107.040 59.380 107.210 ;
        RECT 59.830 107.040 60.170 107.210 ;
        RECT 60.620 107.040 60.960 107.210 ;
        RECT 61.410 107.040 61.750 107.210 ;
        RECT 62.200 107.040 62.540 107.210 ;
        RECT 64.890 107.040 65.230 107.210 ;
        RECT 65.680 107.040 66.020 107.210 ;
        RECT 66.470 107.040 66.810 107.210 ;
        RECT 67.260 107.040 67.600 107.210 ;
        RECT 68.050 107.040 68.390 107.210 ;
        RECT 68.840 107.040 69.180 107.210 ;
        RECT 69.630 107.040 69.970 107.210 ;
        RECT 70.420 107.040 70.760 107.210 ;
        RECT 71.210 107.040 71.550 107.210 ;
        RECT 72.000 107.040 72.340 107.210 ;
        RECT 20.105 106.175 20.445 106.345 ;
        RECT 20.895 106.175 21.235 106.345 ;
        RECT 21.685 106.175 22.025 106.345 ;
        RECT 22.475 106.175 22.815 106.345 ;
        RECT 16.920 103.950 17.260 104.120 ;
        RECT 16.610 102.820 16.780 103.700 ;
        RECT 16.920 102.400 17.260 102.570 ;
        RECT 19.615 101.460 19.955 101.630 ;
        RECT 20.405 101.460 20.745 101.630 ;
        RECT 21.195 101.460 21.535 101.630 ;
        RECT 21.985 101.460 22.325 101.630 ;
        RECT 16.920 100.460 17.260 100.630 ;
        RECT 17.400 96.330 17.570 100.210 ;
        RECT 20.095 96.330 20.265 101.210 ;
        RECT 21.675 96.330 21.845 101.210 ;
        RECT 25.550 96.400 25.890 96.570 ;
        RECT 26.340 96.400 26.680 96.570 ;
        RECT 27.130 96.400 27.470 96.570 ;
        RECT 27.920 96.400 28.260 96.570 ;
        RECT 28.710 96.400 29.050 96.570 ;
        RECT 29.500 96.400 29.840 96.570 ;
        RECT 30.290 96.400 30.630 96.570 ;
        RECT 31.080 96.400 31.420 96.570 ;
        RECT 31.870 96.400 32.210 96.570 ;
        RECT 32.660 96.400 33.000 96.570 ;
        RECT 35.490 96.400 35.830 96.570 ;
        RECT 36.280 96.400 36.620 96.570 ;
        RECT 37.070 96.400 37.410 96.570 ;
        RECT 37.860 96.400 38.200 96.570 ;
        RECT 38.650 96.400 38.990 96.570 ;
        RECT 39.440 96.400 39.780 96.570 ;
        RECT 40.230 96.400 40.570 96.570 ;
        RECT 41.020 96.400 41.360 96.570 ;
        RECT 41.810 96.400 42.150 96.570 ;
        RECT 42.600 96.400 42.940 96.570 ;
        RECT 45.290 96.400 45.630 96.570 ;
        RECT 46.080 96.400 46.420 96.570 ;
        RECT 46.870 96.400 47.210 96.570 ;
        RECT 47.660 96.400 48.000 96.570 ;
        RECT 48.450 96.400 48.790 96.570 ;
        RECT 49.240 96.400 49.580 96.570 ;
        RECT 50.030 96.400 50.370 96.570 ;
        RECT 50.820 96.400 51.160 96.570 ;
        RECT 51.610 96.400 51.950 96.570 ;
        RECT 52.400 96.400 52.740 96.570 ;
        RECT 55.090 96.400 55.430 96.570 ;
        RECT 55.880 96.400 56.220 96.570 ;
        RECT 56.670 96.400 57.010 96.570 ;
        RECT 57.460 96.400 57.800 96.570 ;
        RECT 58.250 96.400 58.590 96.570 ;
        RECT 59.040 96.400 59.380 96.570 ;
        RECT 59.830 96.400 60.170 96.570 ;
        RECT 60.620 96.400 60.960 96.570 ;
        RECT 61.410 96.400 61.750 96.570 ;
        RECT 62.200 96.400 62.540 96.570 ;
        RECT 64.890 96.400 65.230 96.570 ;
        RECT 65.680 96.400 66.020 96.570 ;
        RECT 66.470 96.400 66.810 96.570 ;
        RECT 67.260 96.400 67.600 96.570 ;
        RECT 68.050 96.400 68.390 96.570 ;
        RECT 68.840 96.400 69.180 96.570 ;
        RECT 69.630 96.400 69.970 96.570 ;
        RECT 70.420 96.400 70.760 96.570 ;
        RECT 71.210 96.400 71.550 96.570 ;
        RECT 72.000 96.400 72.340 96.570 ;
        RECT 16.920 95.910 17.260 96.080 ;
        RECT 19.615 95.910 19.955 96.080 ;
        RECT 20.405 95.910 20.745 96.080 ;
        RECT 21.195 95.910 21.535 96.080 ;
        RECT 21.985 95.910 22.325 96.080 ;
        RECT 15.365 93.950 15.705 94.120 ;
        RECT 16.155 93.950 16.495 94.120 ;
        RECT 16.945 93.950 17.285 94.120 ;
        RECT 17.735 93.950 18.075 94.120 ;
        RECT 18.525 93.950 18.865 94.120 ;
        RECT 19.315 93.950 19.655 94.120 ;
        RECT 20.105 93.950 20.445 94.120 ;
        RECT 20.895 93.950 21.235 94.120 ;
        RECT 21.685 93.950 22.025 94.120 ;
        RECT 22.475 93.950 22.815 94.120 ;
        RECT 25.555 93.965 25.895 94.135 ;
        RECT 26.345 93.965 26.685 94.135 ;
        RECT 27.135 93.965 27.475 94.135 ;
        RECT 27.925 93.965 28.265 94.135 ;
        RECT 28.715 93.965 29.055 94.135 ;
        RECT 29.505 93.965 29.845 94.135 ;
        RECT 30.295 93.965 30.635 94.135 ;
        RECT 31.085 93.965 31.425 94.135 ;
        RECT 31.875 93.965 32.215 94.135 ;
        RECT 32.665 93.965 33.005 94.135 ;
        RECT 35.495 93.965 35.835 94.135 ;
        RECT 36.285 93.965 36.625 94.135 ;
        RECT 37.075 93.965 37.415 94.135 ;
        RECT 37.865 93.965 38.205 94.135 ;
        RECT 38.655 93.965 38.995 94.135 ;
        RECT 39.445 93.965 39.785 94.135 ;
        RECT 40.235 93.965 40.575 94.135 ;
        RECT 41.025 93.965 41.365 94.135 ;
        RECT 41.815 93.965 42.155 94.135 ;
        RECT 42.605 93.965 42.945 94.135 ;
        RECT 45.295 93.965 45.635 94.135 ;
        RECT 46.085 93.965 46.425 94.135 ;
        RECT 46.875 93.965 47.215 94.135 ;
        RECT 47.665 93.965 48.005 94.135 ;
        RECT 48.455 93.965 48.795 94.135 ;
        RECT 49.245 93.965 49.585 94.135 ;
        RECT 50.035 93.965 50.375 94.135 ;
        RECT 50.825 93.965 51.165 94.135 ;
        RECT 51.615 93.965 51.955 94.135 ;
        RECT 52.405 93.965 52.745 94.135 ;
        RECT 55.095 93.965 55.435 94.135 ;
        RECT 55.885 93.965 56.225 94.135 ;
        RECT 56.675 93.965 57.015 94.135 ;
        RECT 57.465 93.965 57.805 94.135 ;
        RECT 58.255 93.965 58.595 94.135 ;
        RECT 59.045 93.965 59.385 94.135 ;
        RECT 59.835 93.965 60.175 94.135 ;
        RECT 60.625 93.965 60.965 94.135 ;
        RECT 61.415 93.965 61.755 94.135 ;
        RECT 62.205 93.965 62.545 94.135 ;
        RECT 64.895 93.965 65.235 94.135 ;
        RECT 65.685 93.965 66.025 94.135 ;
        RECT 66.475 93.965 66.815 94.135 ;
        RECT 67.265 93.965 67.605 94.135 ;
        RECT 68.055 93.965 68.395 94.135 ;
        RECT 68.845 93.965 69.185 94.135 ;
        RECT 69.635 93.965 69.975 94.135 ;
        RECT 70.425 93.965 70.765 94.135 ;
        RECT 71.215 93.965 71.555 94.135 ;
        RECT 72.005 93.965 72.345 94.135 ;
        RECT 15.845 83.820 16.015 93.700 ;
        RECT 17.425 83.820 17.595 93.700 ;
        RECT 19.005 83.820 19.175 93.700 ;
        RECT 20.585 83.820 20.755 93.700 ;
        RECT 22.165 83.820 22.335 93.700 ;
        RECT 15.365 83.400 15.705 83.570 ;
        RECT 16.155 83.400 16.495 83.570 ;
        RECT 16.945 83.400 17.285 83.570 ;
        RECT 17.735 83.400 18.075 83.570 ;
        RECT 18.525 83.400 18.865 83.570 ;
        RECT 19.315 83.400 19.655 83.570 ;
        RECT 20.105 83.400 20.445 83.570 ;
        RECT 20.895 83.400 21.235 83.570 ;
        RECT 21.685 83.400 22.025 83.570 ;
        RECT 22.475 83.400 22.815 83.570 ;
        RECT 25.555 83.415 25.895 83.585 ;
        RECT 26.345 83.415 26.685 83.585 ;
        RECT 27.135 83.415 27.475 83.585 ;
        RECT 27.925 83.415 28.265 83.585 ;
        RECT 28.715 83.415 29.055 83.585 ;
        RECT 29.505 83.415 29.845 83.585 ;
        RECT 30.295 83.415 30.635 83.585 ;
        RECT 31.085 83.415 31.425 83.585 ;
        RECT 31.875 83.415 32.215 83.585 ;
        RECT 32.665 83.415 33.005 83.585 ;
        RECT 35.495 83.415 35.835 83.585 ;
        RECT 36.285 83.415 36.625 83.585 ;
        RECT 37.075 83.415 37.415 83.585 ;
        RECT 37.865 83.415 38.205 83.585 ;
        RECT 38.655 83.415 38.995 83.585 ;
        RECT 39.445 83.415 39.785 83.585 ;
        RECT 40.235 83.415 40.575 83.585 ;
        RECT 41.025 83.415 41.365 83.585 ;
        RECT 41.815 83.415 42.155 83.585 ;
        RECT 42.605 83.415 42.945 83.585 ;
        RECT 45.295 83.415 45.635 83.585 ;
        RECT 46.085 83.415 46.425 83.585 ;
        RECT 46.875 83.415 47.215 83.585 ;
        RECT 47.665 83.415 48.005 83.585 ;
        RECT 48.455 83.415 48.795 83.585 ;
        RECT 49.245 83.415 49.585 83.585 ;
        RECT 50.035 83.415 50.375 83.585 ;
        RECT 50.825 83.415 51.165 83.585 ;
        RECT 51.615 83.415 51.955 83.585 ;
        RECT 52.405 83.415 52.745 83.585 ;
        RECT 55.095 83.415 55.435 83.585 ;
        RECT 55.885 83.415 56.225 83.585 ;
        RECT 56.675 83.415 57.015 83.585 ;
        RECT 57.465 83.415 57.805 83.585 ;
        RECT 58.255 83.415 58.595 83.585 ;
        RECT 59.045 83.415 59.385 83.585 ;
        RECT 59.835 83.415 60.175 83.585 ;
        RECT 60.625 83.415 60.965 83.585 ;
        RECT 61.415 83.415 61.755 83.585 ;
        RECT 62.205 83.415 62.545 83.585 ;
        RECT 64.895 83.415 65.235 83.585 ;
        RECT 65.685 83.415 66.025 83.585 ;
        RECT 66.475 83.415 66.815 83.585 ;
        RECT 67.265 83.415 67.605 83.585 ;
        RECT 68.055 83.415 68.395 83.585 ;
        RECT 68.845 83.415 69.185 83.585 ;
        RECT 69.635 83.415 69.975 83.585 ;
        RECT 70.425 83.415 70.765 83.585 ;
        RECT 71.215 83.415 71.555 83.585 ;
        RECT 72.005 83.415 72.345 83.585 ;
        RECT 25.555 82.885 25.895 83.055 ;
        RECT 26.345 82.885 26.685 83.055 ;
        RECT 27.135 82.885 27.475 83.055 ;
        RECT 27.925 82.885 28.265 83.055 ;
        RECT 28.715 82.885 29.055 83.055 ;
        RECT 29.505 82.885 29.845 83.055 ;
        RECT 30.295 82.885 30.635 83.055 ;
        RECT 31.085 82.885 31.425 83.055 ;
        RECT 31.875 82.885 32.215 83.055 ;
        RECT 32.665 82.885 33.005 83.055 ;
        RECT 35.495 82.885 35.835 83.055 ;
        RECT 36.285 82.885 36.625 83.055 ;
        RECT 37.075 82.885 37.415 83.055 ;
        RECT 37.865 82.885 38.205 83.055 ;
        RECT 38.655 82.885 38.995 83.055 ;
        RECT 39.445 82.885 39.785 83.055 ;
        RECT 40.235 82.885 40.575 83.055 ;
        RECT 41.025 82.885 41.365 83.055 ;
        RECT 41.815 82.885 42.155 83.055 ;
        RECT 42.605 82.885 42.945 83.055 ;
        RECT 45.295 82.885 45.635 83.055 ;
        RECT 46.085 82.885 46.425 83.055 ;
        RECT 46.875 82.885 47.215 83.055 ;
        RECT 47.665 82.885 48.005 83.055 ;
        RECT 48.455 82.885 48.795 83.055 ;
        RECT 49.245 82.885 49.585 83.055 ;
        RECT 50.035 82.885 50.375 83.055 ;
        RECT 50.825 82.885 51.165 83.055 ;
        RECT 51.615 82.885 51.955 83.055 ;
        RECT 52.405 82.885 52.745 83.055 ;
        RECT 55.095 82.885 55.435 83.055 ;
        RECT 55.885 82.885 56.225 83.055 ;
        RECT 56.675 82.885 57.015 83.055 ;
        RECT 57.465 82.885 57.805 83.055 ;
        RECT 58.255 82.885 58.595 83.055 ;
        RECT 59.045 82.885 59.385 83.055 ;
        RECT 59.835 82.885 60.175 83.055 ;
        RECT 60.625 82.885 60.965 83.055 ;
        RECT 61.415 82.885 61.755 83.055 ;
        RECT 62.205 82.885 62.545 83.055 ;
        RECT 64.895 82.885 65.235 83.055 ;
        RECT 65.685 82.885 66.025 83.055 ;
        RECT 66.475 82.885 66.815 83.055 ;
        RECT 67.265 82.885 67.605 83.055 ;
        RECT 68.055 82.885 68.395 83.055 ;
        RECT 68.845 82.885 69.185 83.055 ;
        RECT 69.635 82.885 69.975 83.055 ;
        RECT 70.425 82.885 70.765 83.055 ;
        RECT 71.215 82.885 71.555 83.055 ;
        RECT 72.005 82.885 72.345 83.055 ;
        RECT 3.675 80.690 4.015 80.860 ;
        RECT 4.465 80.690 4.805 80.860 ;
        RECT 5.255 80.690 5.595 80.860 ;
        RECT 6.045 80.690 6.385 80.860 ;
        RECT 6.835 80.690 7.175 80.860 ;
        RECT 8.965 80.690 9.305 80.860 ;
        RECT 9.755 80.690 10.095 80.860 ;
        RECT 10.545 80.690 10.885 80.860 ;
        RECT 11.335 80.690 11.675 80.860 ;
        RECT 12.125 80.690 12.465 80.860 ;
        RECT 4.155 78.510 4.325 80.390 ;
        RECT 5.735 78.510 5.905 80.390 ;
        RECT 7.315 78.510 7.485 80.390 ;
        RECT 8.655 78.510 8.825 80.390 ;
        RECT 10.235 78.510 10.405 80.390 ;
        RECT 11.815 78.510 11.985 80.390 ;
        RECT 18.045 80.110 18.385 80.280 ;
        RECT 18.835 80.110 19.175 80.280 ;
        RECT 21.125 80.110 21.465 80.280 ;
        RECT 21.915 80.110 22.255 80.280 ;
        RECT 3.675 78.040 4.015 78.210 ;
        RECT 4.465 78.040 4.805 78.210 ;
        RECT 5.255 78.040 5.595 78.210 ;
        RECT 6.045 78.040 6.385 78.210 ;
        RECT 6.835 78.040 7.175 78.210 ;
        RECT 8.965 78.040 9.305 78.210 ;
        RECT 9.755 78.040 10.095 78.210 ;
        RECT 10.545 78.040 10.885 78.210 ;
        RECT 11.335 78.040 11.675 78.210 ;
        RECT 12.125 78.040 12.465 78.210 ;
        RECT 1.015 65.375 1.185 75.255 ;
        RECT 2.205 65.375 2.375 75.255 ;
        RECT 3.395 65.375 3.565 75.255 ;
        RECT 4.585 65.375 4.755 75.255 ;
        RECT 5.775 65.375 5.945 75.255 ;
        RECT 6.965 65.375 7.135 75.255 ;
        RECT 8.865 65.375 9.035 75.255 ;
        RECT 10.055 65.375 10.225 75.255 ;
        RECT 11.245 65.375 11.415 75.255 ;
        RECT 12.435 65.375 12.605 75.255 ;
        RECT 13.625 65.375 13.795 75.255 ;
        RECT 14.815 65.375 14.985 75.255 ;
        RECT 18.525 69.930 18.695 79.810 ;
        RECT 21.605 69.930 21.775 79.810 ;
        RECT 25.555 72.335 25.895 72.505 ;
        RECT 26.345 72.335 26.685 72.505 ;
        RECT 27.135 72.335 27.475 72.505 ;
        RECT 27.925 72.335 28.265 72.505 ;
        RECT 28.715 72.335 29.055 72.505 ;
        RECT 29.505 72.335 29.845 72.505 ;
        RECT 30.295 72.335 30.635 72.505 ;
        RECT 31.085 72.335 31.425 72.505 ;
        RECT 31.875 72.335 32.215 72.505 ;
        RECT 32.665 72.335 33.005 72.505 ;
        RECT 35.495 72.335 35.835 72.505 ;
        RECT 36.285 72.335 36.625 72.505 ;
        RECT 37.075 72.335 37.415 72.505 ;
        RECT 37.865 72.335 38.205 72.505 ;
        RECT 38.655 72.335 38.995 72.505 ;
        RECT 39.445 72.335 39.785 72.505 ;
        RECT 40.235 72.335 40.575 72.505 ;
        RECT 41.025 72.335 41.365 72.505 ;
        RECT 41.815 72.335 42.155 72.505 ;
        RECT 42.605 72.335 42.945 72.505 ;
        RECT 45.295 72.335 45.635 72.505 ;
        RECT 46.085 72.335 46.425 72.505 ;
        RECT 46.875 72.335 47.215 72.505 ;
        RECT 47.665 72.335 48.005 72.505 ;
        RECT 48.455 72.335 48.795 72.505 ;
        RECT 49.245 72.335 49.585 72.505 ;
        RECT 50.035 72.335 50.375 72.505 ;
        RECT 50.825 72.335 51.165 72.505 ;
        RECT 51.615 72.335 51.955 72.505 ;
        RECT 52.405 72.335 52.745 72.505 ;
        RECT 55.095 72.335 55.435 72.505 ;
        RECT 55.885 72.335 56.225 72.505 ;
        RECT 56.675 72.335 57.015 72.505 ;
        RECT 57.465 72.335 57.805 72.505 ;
        RECT 58.255 72.335 58.595 72.505 ;
        RECT 59.045 72.335 59.385 72.505 ;
        RECT 59.835 72.335 60.175 72.505 ;
        RECT 60.625 72.335 60.965 72.505 ;
        RECT 61.415 72.335 61.755 72.505 ;
        RECT 62.205 72.335 62.545 72.505 ;
        RECT 64.895 72.335 65.235 72.505 ;
        RECT 65.685 72.335 66.025 72.505 ;
        RECT 66.475 72.335 66.815 72.505 ;
        RECT 67.265 72.335 67.605 72.505 ;
        RECT 68.055 72.335 68.395 72.505 ;
        RECT 68.845 72.335 69.185 72.505 ;
        RECT 69.635 72.335 69.975 72.505 ;
        RECT 70.425 72.335 70.765 72.505 ;
        RECT 71.215 72.335 71.555 72.505 ;
        RECT 72.005 72.335 72.345 72.505 ;
        RECT 18.045 69.460 18.385 69.630 ;
        RECT 18.835 69.460 19.175 69.630 ;
        RECT 21.125 69.460 21.465 69.630 ;
        RECT 21.915 69.460 22.255 69.630 ;
        RECT 25.555 69.325 25.895 69.495 ;
        RECT 26.345 69.325 26.685 69.495 ;
        RECT 27.135 69.325 27.475 69.495 ;
        RECT 27.925 69.325 28.265 69.495 ;
        RECT 28.715 69.325 29.055 69.495 ;
        RECT 29.505 69.325 29.845 69.495 ;
        RECT 30.295 69.325 30.635 69.495 ;
        RECT 31.085 69.325 31.425 69.495 ;
        RECT 31.875 69.325 32.215 69.495 ;
        RECT 32.665 69.325 33.005 69.495 ;
        RECT 35.495 69.325 35.835 69.495 ;
        RECT 36.285 69.325 36.625 69.495 ;
        RECT 37.075 69.325 37.415 69.495 ;
        RECT 37.865 69.325 38.205 69.495 ;
        RECT 38.655 69.325 38.995 69.495 ;
        RECT 39.445 69.325 39.785 69.495 ;
        RECT 40.235 69.325 40.575 69.495 ;
        RECT 41.025 69.325 41.365 69.495 ;
        RECT 41.815 69.325 42.155 69.495 ;
        RECT 42.605 69.325 42.945 69.495 ;
        RECT 45.295 69.325 45.635 69.495 ;
        RECT 46.085 69.325 46.425 69.495 ;
        RECT 46.875 69.325 47.215 69.495 ;
        RECT 47.665 69.325 48.005 69.495 ;
        RECT 48.455 69.325 48.795 69.495 ;
        RECT 49.245 69.325 49.585 69.495 ;
        RECT 50.035 69.325 50.375 69.495 ;
        RECT 50.825 69.325 51.165 69.495 ;
        RECT 51.615 69.325 51.955 69.495 ;
        RECT 52.405 69.325 52.745 69.495 ;
        RECT 55.095 69.325 55.435 69.495 ;
        RECT 55.885 69.325 56.225 69.495 ;
        RECT 56.675 69.325 57.015 69.495 ;
        RECT 57.465 69.325 57.805 69.495 ;
        RECT 58.255 69.325 58.595 69.495 ;
        RECT 59.045 69.325 59.385 69.495 ;
        RECT 59.835 69.325 60.175 69.495 ;
        RECT 60.625 69.325 60.965 69.495 ;
        RECT 61.415 69.325 61.755 69.495 ;
        RECT 62.205 69.325 62.545 69.495 ;
        RECT 64.895 69.325 65.235 69.495 ;
        RECT 65.685 69.325 66.025 69.495 ;
        RECT 66.475 69.325 66.815 69.495 ;
        RECT 67.265 69.325 67.605 69.495 ;
        RECT 68.055 69.325 68.395 69.495 ;
        RECT 68.845 69.325 69.185 69.495 ;
        RECT 69.635 69.325 69.975 69.495 ;
        RECT 70.425 69.325 70.765 69.495 ;
        RECT 71.215 69.325 71.555 69.495 ;
        RECT 72.005 69.325 72.345 69.495 ;
        RECT 18.045 67.030 18.385 67.200 ;
        RECT 18.835 67.030 19.175 67.200 ;
        RECT 21.125 67.030 21.465 67.200 ;
        RECT 21.915 67.030 22.255 67.200 ;
        RECT 3.105 60.810 3.275 62.690 ;
        RECT 4.065 60.810 4.235 62.690 ;
        RECT 5.025 60.810 5.195 62.690 ;
        RECT 5.975 60.810 6.145 62.690 ;
        RECT 6.935 60.810 7.105 62.690 ;
        RECT 9.035 60.810 9.205 62.690 ;
        RECT 9.995 60.810 10.165 62.690 ;
        RECT 10.955 60.810 11.125 62.690 ;
        RECT 11.905 60.810 12.075 62.690 ;
        RECT 12.865 60.810 13.035 62.690 ;
        RECT 18.525 61.900 18.695 66.780 ;
        RECT 21.605 61.900 21.775 66.780 ;
        RECT 18.045 61.480 18.385 61.650 ;
        RECT 18.835 61.480 19.175 61.650 ;
        RECT 21.125 61.480 21.465 61.650 ;
        RECT 21.915 61.480 22.255 61.650 ;
        RECT 25.555 58.775 25.895 58.945 ;
        RECT 26.345 58.775 26.685 58.945 ;
        RECT 27.135 58.775 27.475 58.945 ;
        RECT 27.925 58.775 28.265 58.945 ;
        RECT 28.715 58.775 29.055 58.945 ;
        RECT 29.505 58.775 29.845 58.945 ;
        RECT 30.295 58.775 30.635 58.945 ;
        RECT 31.085 58.775 31.425 58.945 ;
        RECT 31.875 58.775 32.215 58.945 ;
        RECT 32.665 58.775 33.005 58.945 ;
        RECT 35.495 58.775 35.835 58.945 ;
        RECT 36.285 58.775 36.625 58.945 ;
        RECT 37.075 58.775 37.415 58.945 ;
        RECT 37.865 58.775 38.205 58.945 ;
        RECT 38.655 58.775 38.995 58.945 ;
        RECT 39.445 58.775 39.785 58.945 ;
        RECT 40.235 58.775 40.575 58.945 ;
        RECT 41.025 58.775 41.365 58.945 ;
        RECT 41.815 58.775 42.155 58.945 ;
        RECT 42.605 58.775 42.945 58.945 ;
        RECT 45.295 58.775 45.635 58.945 ;
        RECT 46.085 58.775 46.425 58.945 ;
        RECT 46.875 58.775 47.215 58.945 ;
        RECT 47.665 58.775 48.005 58.945 ;
        RECT 48.455 58.775 48.795 58.945 ;
        RECT 49.245 58.775 49.585 58.945 ;
        RECT 50.035 58.775 50.375 58.945 ;
        RECT 50.825 58.775 51.165 58.945 ;
        RECT 51.615 58.775 51.955 58.945 ;
        RECT 52.405 58.775 52.745 58.945 ;
        RECT 55.095 58.775 55.435 58.945 ;
        RECT 55.885 58.775 56.225 58.945 ;
        RECT 56.675 58.775 57.015 58.945 ;
        RECT 57.465 58.775 57.805 58.945 ;
        RECT 58.255 58.775 58.595 58.945 ;
        RECT 59.045 58.775 59.385 58.945 ;
        RECT 59.835 58.775 60.175 58.945 ;
        RECT 60.625 58.775 60.965 58.945 ;
        RECT 61.415 58.775 61.755 58.945 ;
        RECT 62.205 58.775 62.545 58.945 ;
        RECT 64.895 58.775 65.235 58.945 ;
        RECT 65.685 58.775 66.025 58.945 ;
        RECT 66.475 58.775 66.815 58.945 ;
        RECT 67.265 58.775 67.605 58.945 ;
        RECT 68.055 58.775 68.395 58.945 ;
        RECT 68.845 58.775 69.185 58.945 ;
        RECT 69.635 58.775 69.975 58.945 ;
        RECT 70.425 58.775 70.765 58.945 ;
        RECT 71.215 58.775 71.555 58.945 ;
        RECT 72.005 58.775 72.345 58.945 ;
        RECT 15.365 58.260 15.705 58.430 ;
        RECT 16.155 58.260 16.495 58.430 ;
        RECT 16.945 58.260 17.285 58.430 ;
        RECT 17.735 58.260 18.075 58.430 ;
        RECT 18.525 58.260 18.865 58.430 ;
        RECT 19.315 58.260 19.655 58.430 ;
        RECT 20.105 58.260 20.445 58.430 ;
        RECT 20.895 58.260 21.235 58.430 ;
        RECT 21.685 58.260 22.025 58.430 ;
        RECT 22.475 58.260 22.815 58.430 ;
        RECT 25.555 58.245 25.895 58.415 ;
        RECT 26.345 58.245 26.685 58.415 ;
        RECT 27.135 58.245 27.475 58.415 ;
        RECT 27.925 58.245 28.265 58.415 ;
        RECT 28.715 58.245 29.055 58.415 ;
        RECT 29.505 58.245 29.845 58.415 ;
        RECT 30.295 58.245 30.635 58.415 ;
        RECT 31.085 58.245 31.425 58.415 ;
        RECT 31.875 58.245 32.215 58.415 ;
        RECT 32.665 58.245 33.005 58.415 ;
        RECT 35.495 58.245 35.835 58.415 ;
        RECT 36.285 58.245 36.625 58.415 ;
        RECT 37.075 58.245 37.415 58.415 ;
        RECT 37.865 58.245 38.205 58.415 ;
        RECT 38.655 58.245 38.995 58.415 ;
        RECT 39.445 58.245 39.785 58.415 ;
        RECT 40.235 58.245 40.575 58.415 ;
        RECT 41.025 58.245 41.365 58.415 ;
        RECT 41.815 58.245 42.155 58.415 ;
        RECT 42.605 58.245 42.945 58.415 ;
        RECT 45.295 58.245 45.635 58.415 ;
        RECT 46.085 58.245 46.425 58.415 ;
        RECT 46.875 58.245 47.215 58.415 ;
        RECT 47.665 58.245 48.005 58.415 ;
        RECT 48.455 58.245 48.795 58.415 ;
        RECT 49.245 58.245 49.585 58.415 ;
        RECT 50.035 58.245 50.375 58.415 ;
        RECT 50.825 58.245 51.165 58.415 ;
        RECT 51.615 58.245 51.955 58.415 ;
        RECT 52.405 58.245 52.745 58.415 ;
        RECT 55.095 58.245 55.435 58.415 ;
        RECT 55.885 58.245 56.225 58.415 ;
        RECT 56.675 58.245 57.015 58.415 ;
        RECT 57.465 58.245 57.805 58.415 ;
        RECT 58.255 58.245 58.595 58.415 ;
        RECT 59.045 58.245 59.385 58.415 ;
        RECT 59.835 58.245 60.175 58.415 ;
        RECT 60.625 58.245 60.965 58.415 ;
        RECT 61.415 58.245 61.755 58.415 ;
        RECT 62.205 58.245 62.545 58.415 ;
        RECT 64.895 58.245 65.235 58.415 ;
        RECT 65.685 58.245 66.025 58.415 ;
        RECT 66.475 58.245 66.815 58.415 ;
        RECT 67.265 58.245 67.605 58.415 ;
        RECT 68.055 58.245 68.395 58.415 ;
        RECT 68.845 58.245 69.185 58.415 ;
        RECT 69.635 58.245 69.975 58.415 ;
        RECT 70.425 58.245 70.765 58.415 ;
        RECT 71.215 58.245 71.555 58.415 ;
        RECT 72.005 58.245 72.345 58.415 ;
        RECT 15.845 48.130 16.015 58.010 ;
        RECT 17.425 48.130 17.595 58.010 ;
        RECT 19.005 48.130 19.175 58.010 ;
        RECT 20.585 48.130 20.755 58.010 ;
        RECT 22.165 48.130 22.335 58.010 ;
        RECT 15.365 47.710 15.705 47.880 ;
        RECT 16.155 47.710 16.495 47.880 ;
        RECT 16.945 47.710 17.285 47.880 ;
        RECT 17.735 47.710 18.075 47.880 ;
        RECT 18.525 47.710 18.865 47.880 ;
        RECT 19.315 47.710 19.655 47.880 ;
        RECT 20.105 47.710 20.445 47.880 ;
        RECT 20.895 47.710 21.235 47.880 ;
        RECT 21.685 47.710 22.025 47.880 ;
        RECT 22.475 47.710 22.815 47.880 ;
        RECT 25.555 47.695 25.895 47.865 ;
        RECT 26.345 47.695 26.685 47.865 ;
        RECT 27.135 47.695 27.475 47.865 ;
        RECT 27.925 47.695 28.265 47.865 ;
        RECT 28.715 47.695 29.055 47.865 ;
        RECT 29.505 47.695 29.845 47.865 ;
        RECT 30.295 47.695 30.635 47.865 ;
        RECT 31.085 47.695 31.425 47.865 ;
        RECT 31.875 47.695 32.215 47.865 ;
        RECT 32.665 47.695 33.005 47.865 ;
        RECT 35.495 47.695 35.835 47.865 ;
        RECT 36.285 47.695 36.625 47.865 ;
        RECT 37.075 47.695 37.415 47.865 ;
        RECT 37.865 47.695 38.205 47.865 ;
        RECT 38.655 47.695 38.995 47.865 ;
        RECT 39.445 47.695 39.785 47.865 ;
        RECT 40.235 47.695 40.575 47.865 ;
        RECT 41.025 47.695 41.365 47.865 ;
        RECT 41.815 47.695 42.155 47.865 ;
        RECT 42.605 47.695 42.945 47.865 ;
        RECT 45.295 47.695 45.635 47.865 ;
        RECT 46.085 47.695 46.425 47.865 ;
        RECT 46.875 47.695 47.215 47.865 ;
        RECT 47.665 47.695 48.005 47.865 ;
        RECT 48.455 47.695 48.795 47.865 ;
        RECT 49.245 47.695 49.585 47.865 ;
        RECT 50.035 47.695 50.375 47.865 ;
        RECT 50.825 47.695 51.165 47.865 ;
        RECT 51.615 47.695 51.955 47.865 ;
        RECT 52.405 47.695 52.745 47.865 ;
        RECT 55.095 47.695 55.435 47.865 ;
        RECT 55.885 47.695 56.225 47.865 ;
        RECT 56.675 47.695 57.015 47.865 ;
        RECT 57.465 47.695 57.805 47.865 ;
        RECT 58.255 47.695 58.595 47.865 ;
        RECT 59.045 47.695 59.385 47.865 ;
        RECT 59.835 47.695 60.175 47.865 ;
        RECT 60.625 47.695 60.965 47.865 ;
        RECT 61.415 47.695 61.755 47.865 ;
        RECT 62.205 47.695 62.545 47.865 ;
        RECT 64.895 47.695 65.235 47.865 ;
        RECT 65.685 47.695 66.025 47.865 ;
        RECT 66.475 47.695 66.815 47.865 ;
        RECT 67.265 47.695 67.605 47.865 ;
        RECT 68.055 47.695 68.395 47.865 ;
        RECT 68.845 47.695 69.185 47.865 ;
        RECT 69.635 47.695 69.975 47.865 ;
        RECT 70.425 47.695 70.765 47.865 ;
        RECT 71.215 47.695 71.555 47.865 ;
        RECT 72.005 47.695 72.345 47.865 ;
        RECT 16.920 45.750 17.260 45.920 ;
        RECT 19.615 45.750 19.955 45.920 ;
        RECT 20.405 45.750 20.745 45.920 ;
        RECT 21.195 45.750 21.535 45.920 ;
        RECT 21.985 45.750 22.325 45.920 ;
        RECT 17.400 41.620 17.570 45.500 ;
        RECT 16.920 41.200 17.260 41.370 ;
        RECT 20.095 40.620 20.265 45.500 ;
        RECT 21.675 40.620 21.845 45.500 ;
        RECT 25.550 45.260 25.890 45.430 ;
        RECT 26.340 45.260 26.680 45.430 ;
        RECT 27.130 45.260 27.470 45.430 ;
        RECT 27.920 45.260 28.260 45.430 ;
        RECT 28.710 45.260 29.050 45.430 ;
        RECT 29.500 45.260 29.840 45.430 ;
        RECT 30.290 45.260 30.630 45.430 ;
        RECT 31.080 45.260 31.420 45.430 ;
        RECT 31.870 45.260 32.210 45.430 ;
        RECT 32.660 45.260 33.000 45.430 ;
        RECT 35.490 45.260 35.830 45.430 ;
        RECT 36.280 45.260 36.620 45.430 ;
        RECT 37.070 45.260 37.410 45.430 ;
        RECT 37.860 45.260 38.200 45.430 ;
        RECT 38.650 45.260 38.990 45.430 ;
        RECT 39.440 45.260 39.780 45.430 ;
        RECT 40.230 45.260 40.570 45.430 ;
        RECT 41.020 45.260 41.360 45.430 ;
        RECT 41.810 45.260 42.150 45.430 ;
        RECT 42.600 45.260 42.940 45.430 ;
        RECT 45.290 45.260 45.630 45.430 ;
        RECT 46.080 45.260 46.420 45.430 ;
        RECT 46.870 45.260 47.210 45.430 ;
        RECT 47.660 45.260 48.000 45.430 ;
        RECT 48.450 45.260 48.790 45.430 ;
        RECT 49.240 45.260 49.580 45.430 ;
        RECT 50.030 45.260 50.370 45.430 ;
        RECT 50.820 45.260 51.160 45.430 ;
        RECT 51.610 45.260 51.950 45.430 ;
        RECT 52.400 45.260 52.740 45.430 ;
        RECT 55.090 45.260 55.430 45.430 ;
        RECT 55.880 45.260 56.220 45.430 ;
        RECT 56.670 45.260 57.010 45.430 ;
        RECT 57.460 45.260 57.800 45.430 ;
        RECT 58.250 45.260 58.590 45.430 ;
        RECT 59.040 45.260 59.380 45.430 ;
        RECT 59.830 45.260 60.170 45.430 ;
        RECT 60.620 45.260 60.960 45.430 ;
        RECT 61.410 45.260 61.750 45.430 ;
        RECT 62.200 45.260 62.540 45.430 ;
        RECT 64.890 45.260 65.230 45.430 ;
        RECT 65.680 45.260 66.020 45.430 ;
        RECT 66.470 45.260 66.810 45.430 ;
        RECT 67.260 45.260 67.600 45.430 ;
        RECT 68.050 45.260 68.390 45.430 ;
        RECT 68.840 45.260 69.180 45.430 ;
        RECT 69.630 45.260 69.970 45.430 ;
        RECT 70.420 45.260 70.760 45.430 ;
        RECT 71.210 45.260 71.550 45.430 ;
        RECT 72.000 45.260 72.340 45.430 ;
        RECT 19.615 40.200 19.955 40.370 ;
        RECT 20.405 40.200 20.745 40.370 ;
        RECT 21.195 40.200 21.535 40.370 ;
        RECT 21.985 40.200 22.325 40.370 ;
        RECT 16.920 39.260 17.260 39.430 ;
        RECT 16.610 38.130 16.780 39.010 ;
        RECT 16.920 37.710 17.260 37.880 ;
        RECT 20.105 35.485 20.445 35.655 ;
        RECT 20.895 35.485 21.235 35.655 ;
        RECT 21.685 35.485 22.025 35.655 ;
        RECT 22.475 35.485 22.815 35.655 ;
        RECT 16.615 33.050 16.955 33.220 ;
        RECT 17.405 33.050 17.745 33.220 ;
        RECT 16.305 31.870 16.475 32.750 ;
        RECT 17.885 31.870 18.055 32.750 ;
        RECT 16.620 29.490 16.960 29.660 ;
        RECT 17.410 29.490 17.750 29.660 ;
        RECT 17.100 25.310 17.270 29.190 ;
        RECT 20.585 25.305 20.755 35.185 ;
        RECT 22.165 25.305 22.335 35.185 ;
        RECT 25.550 34.620 25.890 34.790 ;
        RECT 26.340 34.620 26.680 34.790 ;
        RECT 27.130 34.620 27.470 34.790 ;
        RECT 27.920 34.620 28.260 34.790 ;
        RECT 28.710 34.620 29.050 34.790 ;
        RECT 29.500 34.620 29.840 34.790 ;
        RECT 30.290 34.620 30.630 34.790 ;
        RECT 31.080 34.620 31.420 34.790 ;
        RECT 31.870 34.620 32.210 34.790 ;
        RECT 32.660 34.620 33.000 34.790 ;
        RECT 35.490 34.620 35.830 34.790 ;
        RECT 36.280 34.620 36.620 34.790 ;
        RECT 37.070 34.620 37.410 34.790 ;
        RECT 37.860 34.620 38.200 34.790 ;
        RECT 38.650 34.620 38.990 34.790 ;
        RECT 39.440 34.620 39.780 34.790 ;
        RECT 40.230 34.620 40.570 34.790 ;
        RECT 41.020 34.620 41.360 34.790 ;
        RECT 41.810 34.620 42.150 34.790 ;
        RECT 42.600 34.620 42.940 34.790 ;
        RECT 45.290 34.620 45.630 34.790 ;
        RECT 46.080 34.620 46.420 34.790 ;
        RECT 46.870 34.620 47.210 34.790 ;
        RECT 47.660 34.620 48.000 34.790 ;
        RECT 48.450 34.620 48.790 34.790 ;
        RECT 49.240 34.620 49.580 34.790 ;
        RECT 50.030 34.620 50.370 34.790 ;
        RECT 50.820 34.620 51.160 34.790 ;
        RECT 51.610 34.620 51.950 34.790 ;
        RECT 52.400 34.620 52.740 34.790 ;
        RECT 55.090 34.620 55.430 34.790 ;
        RECT 55.880 34.620 56.220 34.790 ;
        RECT 56.670 34.620 57.010 34.790 ;
        RECT 57.460 34.620 57.800 34.790 ;
        RECT 58.250 34.620 58.590 34.790 ;
        RECT 59.040 34.620 59.380 34.790 ;
        RECT 59.830 34.620 60.170 34.790 ;
        RECT 60.620 34.620 60.960 34.790 ;
        RECT 61.410 34.620 61.750 34.790 ;
        RECT 62.200 34.620 62.540 34.790 ;
        RECT 64.890 34.620 65.230 34.790 ;
        RECT 65.680 34.620 66.020 34.790 ;
        RECT 66.470 34.620 66.810 34.790 ;
        RECT 67.260 34.620 67.600 34.790 ;
        RECT 68.050 34.620 68.390 34.790 ;
        RECT 68.840 34.620 69.180 34.790 ;
        RECT 69.630 34.620 69.970 34.790 ;
        RECT 70.420 34.620 70.760 34.790 ;
        RECT 71.210 34.620 71.550 34.790 ;
        RECT 72.000 34.620 72.340 34.790 ;
        RECT 25.550 34.080 25.890 34.250 ;
        RECT 26.340 34.080 26.680 34.250 ;
        RECT 27.130 34.080 27.470 34.250 ;
        RECT 27.920 34.080 28.260 34.250 ;
        RECT 28.710 34.080 29.050 34.250 ;
        RECT 29.500 34.080 29.840 34.250 ;
        RECT 30.290 34.080 30.630 34.250 ;
        RECT 31.080 34.080 31.420 34.250 ;
        RECT 31.870 34.080 32.210 34.250 ;
        RECT 32.660 34.080 33.000 34.250 ;
        RECT 35.490 34.080 35.830 34.250 ;
        RECT 36.280 34.080 36.620 34.250 ;
        RECT 37.070 34.080 37.410 34.250 ;
        RECT 37.860 34.080 38.200 34.250 ;
        RECT 38.650 34.080 38.990 34.250 ;
        RECT 39.440 34.080 39.780 34.250 ;
        RECT 40.230 34.080 40.570 34.250 ;
        RECT 41.020 34.080 41.360 34.250 ;
        RECT 41.810 34.080 42.150 34.250 ;
        RECT 42.600 34.080 42.940 34.250 ;
        RECT 45.290 34.080 45.630 34.250 ;
        RECT 46.080 34.080 46.420 34.250 ;
        RECT 46.870 34.080 47.210 34.250 ;
        RECT 47.660 34.080 48.000 34.250 ;
        RECT 48.450 34.080 48.790 34.250 ;
        RECT 49.240 34.080 49.580 34.250 ;
        RECT 50.030 34.080 50.370 34.250 ;
        RECT 50.820 34.080 51.160 34.250 ;
        RECT 51.610 34.080 51.950 34.250 ;
        RECT 52.400 34.080 52.740 34.250 ;
        RECT 55.090 34.080 55.430 34.250 ;
        RECT 55.880 34.080 56.220 34.250 ;
        RECT 56.670 34.080 57.010 34.250 ;
        RECT 57.460 34.080 57.800 34.250 ;
        RECT 58.250 34.080 58.590 34.250 ;
        RECT 59.040 34.080 59.380 34.250 ;
        RECT 59.830 34.080 60.170 34.250 ;
        RECT 60.620 34.080 60.960 34.250 ;
        RECT 61.410 34.080 61.750 34.250 ;
        RECT 62.200 34.080 62.540 34.250 ;
        RECT 64.890 34.080 65.230 34.250 ;
        RECT 65.680 34.080 66.020 34.250 ;
        RECT 66.470 34.080 66.810 34.250 ;
        RECT 67.260 34.080 67.600 34.250 ;
        RECT 68.050 34.080 68.390 34.250 ;
        RECT 68.840 34.080 69.180 34.250 ;
        RECT 69.630 34.080 69.970 34.250 ;
        RECT 70.420 34.080 70.760 34.250 ;
        RECT 71.210 34.080 71.550 34.250 ;
        RECT 72.000 34.080 72.340 34.250 ;
        RECT 16.620 24.840 16.960 25.010 ;
        RECT 17.410 24.840 17.750 25.010 ;
        RECT 20.105 24.835 20.445 25.005 ;
        RECT 20.895 24.835 21.235 25.005 ;
        RECT 21.685 24.835 22.025 25.005 ;
        RECT 22.475 24.835 22.815 25.005 ;
        RECT 25.550 23.440 25.890 23.610 ;
        RECT 26.340 23.440 26.680 23.610 ;
        RECT 27.130 23.440 27.470 23.610 ;
        RECT 27.920 23.440 28.260 23.610 ;
        RECT 28.710 23.440 29.050 23.610 ;
        RECT 29.500 23.440 29.840 23.610 ;
        RECT 30.290 23.440 30.630 23.610 ;
        RECT 31.080 23.440 31.420 23.610 ;
        RECT 31.870 23.440 32.210 23.610 ;
        RECT 32.660 23.440 33.000 23.610 ;
        RECT 35.490 23.440 35.830 23.610 ;
        RECT 36.280 23.440 36.620 23.610 ;
        RECT 37.070 23.440 37.410 23.610 ;
        RECT 37.860 23.440 38.200 23.610 ;
        RECT 38.650 23.440 38.990 23.610 ;
        RECT 39.440 23.440 39.780 23.610 ;
        RECT 40.230 23.440 40.570 23.610 ;
        RECT 41.020 23.440 41.360 23.610 ;
        RECT 41.810 23.440 42.150 23.610 ;
        RECT 42.600 23.440 42.940 23.610 ;
        RECT 45.290 23.440 45.630 23.610 ;
        RECT 46.080 23.440 46.420 23.610 ;
        RECT 46.870 23.440 47.210 23.610 ;
        RECT 47.660 23.440 48.000 23.610 ;
        RECT 48.450 23.440 48.790 23.610 ;
        RECT 49.240 23.440 49.580 23.610 ;
        RECT 50.030 23.440 50.370 23.610 ;
        RECT 50.820 23.440 51.160 23.610 ;
        RECT 51.610 23.440 51.950 23.610 ;
        RECT 52.400 23.440 52.740 23.610 ;
        RECT 55.090 23.440 55.430 23.610 ;
        RECT 55.880 23.440 56.220 23.610 ;
        RECT 56.670 23.440 57.010 23.610 ;
        RECT 57.460 23.440 57.800 23.610 ;
        RECT 58.250 23.440 58.590 23.610 ;
        RECT 59.040 23.440 59.380 23.610 ;
        RECT 59.830 23.440 60.170 23.610 ;
        RECT 60.620 23.440 60.960 23.610 ;
        RECT 61.410 23.440 61.750 23.610 ;
        RECT 62.200 23.440 62.540 23.610 ;
        RECT 64.890 23.440 65.230 23.610 ;
        RECT 65.680 23.440 66.020 23.610 ;
        RECT 66.470 23.440 66.810 23.610 ;
        RECT 67.260 23.440 67.600 23.610 ;
        RECT 68.050 23.440 68.390 23.610 ;
        RECT 68.840 23.440 69.180 23.610 ;
        RECT 69.630 23.440 69.970 23.610 ;
        RECT 70.420 23.440 70.760 23.610 ;
        RECT 71.210 23.440 71.550 23.610 ;
        RECT 72.000 23.440 72.340 23.610 ;
        RECT 15.365 22.905 15.705 23.075 ;
        RECT 16.155 22.905 16.495 23.075 ;
        RECT 16.945 22.905 17.285 23.075 ;
        RECT 17.735 22.905 18.075 23.075 ;
        RECT 18.525 22.905 18.865 23.075 ;
        RECT 19.315 22.905 19.655 23.075 ;
        RECT 20.105 22.905 20.445 23.075 ;
        RECT 20.895 22.905 21.235 23.075 ;
        RECT 21.685 22.905 22.025 23.075 ;
        RECT 22.475 22.905 22.815 23.075 ;
        RECT 25.550 22.900 25.890 23.070 ;
        RECT 26.340 22.900 26.680 23.070 ;
        RECT 27.130 22.900 27.470 23.070 ;
        RECT 27.920 22.900 28.260 23.070 ;
        RECT 28.710 22.900 29.050 23.070 ;
        RECT 29.500 22.900 29.840 23.070 ;
        RECT 30.290 22.900 30.630 23.070 ;
        RECT 31.080 22.900 31.420 23.070 ;
        RECT 31.870 22.900 32.210 23.070 ;
        RECT 32.660 22.900 33.000 23.070 ;
        RECT 35.490 22.900 35.830 23.070 ;
        RECT 36.280 22.900 36.620 23.070 ;
        RECT 37.070 22.900 37.410 23.070 ;
        RECT 37.860 22.900 38.200 23.070 ;
        RECT 38.650 22.900 38.990 23.070 ;
        RECT 39.440 22.900 39.780 23.070 ;
        RECT 40.230 22.900 40.570 23.070 ;
        RECT 41.020 22.900 41.360 23.070 ;
        RECT 41.810 22.900 42.150 23.070 ;
        RECT 42.600 22.900 42.940 23.070 ;
        RECT 45.290 22.900 45.630 23.070 ;
        RECT 46.080 22.900 46.420 23.070 ;
        RECT 46.870 22.900 47.210 23.070 ;
        RECT 47.660 22.900 48.000 23.070 ;
        RECT 48.450 22.900 48.790 23.070 ;
        RECT 49.240 22.900 49.580 23.070 ;
        RECT 50.030 22.900 50.370 23.070 ;
        RECT 50.820 22.900 51.160 23.070 ;
        RECT 51.610 22.900 51.950 23.070 ;
        RECT 52.400 22.900 52.740 23.070 ;
        RECT 55.090 22.900 55.430 23.070 ;
        RECT 55.880 22.900 56.220 23.070 ;
        RECT 56.670 22.900 57.010 23.070 ;
        RECT 57.460 22.900 57.800 23.070 ;
        RECT 58.250 22.900 58.590 23.070 ;
        RECT 59.040 22.900 59.380 23.070 ;
        RECT 59.830 22.900 60.170 23.070 ;
        RECT 60.620 22.900 60.960 23.070 ;
        RECT 61.410 22.900 61.750 23.070 ;
        RECT 62.200 22.900 62.540 23.070 ;
        RECT 64.890 22.900 65.230 23.070 ;
        RECT 65.680 22.900 66.020 23.070 ;
        RECT 66.470 22.900 66.810 23.070 ;
        RECT 67.260 22.900 67.600 23.070 ;
        RECT 68.050 22.900 68.390 23.070 ;
        RECT 68.840 22.900 69.180 23.070 ;
        RECT 69.630 22.900 69.970 23.070 ;
        RECT 70.420 22.900 70.760 23.070 ;
        RECT 71.210 22.900 71.550 23.070 ;
        RECT 72.000 22.900 72.340 23.070 ;
        RECT 15.845 12.725 16.015 22.605 ;
        RECT 17.425 12.725 17.595 22.605 ;
        RECT 19.005 12.725 19.175 22.605 ;
        RECT 20.585 12.725 20.755 22.605 ;
        RECT 22.165 12.725 22.335 22.605 ;
        RECT 15.365 12.255 15.705 12.425 ;
        RECT 16.155 12.255 16.495 12.425 ;
        RECT 16.945 12.255 17.285 12.425 ;
        RECT 17.735 12.255 18.075 12.425 ;
        RECT 18.525 12.255 18.865 12.425 ;
        RECT 19.315 12.255 19.655 12.425 ;
        RECT 20.105 12.255 20.445 12.425 ;
        RECT 20.895 12.255 21.235 12.425 ;
        RECT 21.685 12.255 22.025 12.425 ;
        RECT 22.475 12.255 22.815 12.425 ;
        RECT 25.550 12.260 25.890 12.430 ;
        RECT 26.340 12.260 26.680 12.430 ;
        RECT 27.130 12.260 27.470 12.430 ;
        RECT 27.920 12.260 28.260 12.430 ;
        RECT 28.710 12.260 29.050 12.430 ;
        RECT 29.500 12.260 29.840 12.430 ;
        RECT 30.290 12.260 30.630 12.430 ;
        RECT 31.080 12.260 31.420 12.430 ;
        RECT 31.870 12.260 32.210 12.430 ;
        RECT 32.660 12.260 33.000 12.430 ;
        RECT 35.490 12.260 35.830 12.430 ;
        RECT 36.280 12.260 36.620 12.430 ;
        RECT 37.070 12.260 37.410 12.430 ;
        RECT 37.860 12.260 38.200 12.430 ;
        RECT 38.650 12.260 38.990 12.430 ;
        RECT 39.440 12.260 39.780 12.430 ;
        RECT 40.230 12.260 40.570 12.430 ;
        RECT 41.020 12.260 41.360 12.430 ;
        RECT 41.810 12.260 42.150 12.430 ;
        RECT 42.600 12.260 42.940 12.430 ;
        RECT 45.290 12.260 45.630 12.430 ;
        RECT 46.080 12.260 46.420 12.430 ;
        RECT 46.870 12.260 47.210 12.430 ;
        RECT 47.660 12.260 48.000 12.430 ;
        RECT 48.450 12.260 48.790 12.430 ;
        RECT 49.240 12.260 49.580 12.430 ;
        RECT 50.030 12.260 50.370 12.430 ;
        RECT 50.820 12.260 51.160 12.430 ;
        RECT 51.610 12.260 51.950 12.430 ;
        RECT 52.400 12.260 52.740 12.430 ;
        RECT 55.090 12.260 55.430 12.430 ;
        RECT 55.880 12.260 56.220 12.430 ;
        RECT 56.670 12.260 57.010 12.430 ;
        RECT 57.460 12.260 57.800 12.430 ;
        RECT 58.250 12.260 58.590 12.430 ;
        RECT 59.040 12.260 59.380 12.430 ;
        RECT 59.830 12.260 60.170 12.430 ;
        RECT 60.620 12.260 60.960 12.430 ;
        RECT 61.410 12.260 61.750 12.430 ;
        RECT 62.200 12.260 62.540 12.430 ;
        RECT 64.890 12.260 65.230 12.430 ;
        RECT 65.680 12.260 66.020 12.430 ;
        RECT 66.470 12.260 66.810 12.430 ;
        RECT 67.260 12.260 67.600 12.430 ;
        RECT 68.050 12.260 68.390 12.430 ;
        RECT 68.840 12.260 69.180 12.430 ;
        RECT 69.630 12.260 69.970 12.430 ;
        RECT 70.420 12.260 70.760 12.430 ;
        RECT 71.210 12.260 71.550 12.430 ;
        RECT 72.000 12.260 72.340 12.430 ;
        RECT 15.365 11.725 15.705 11.895 ;
        RECT 16.155 11.725 16.495 11.895 ;
        RECT 16.945 11.725 17.285 11.895 ;
        RECT 17.735 11.725 18.075 11.895 ;
        RECT 18.525 11.725 18.865 11.895 ;
        RECT 19.315 11.725 19.655 11.895 ;
        RECT 20.105 11.725 20.445 11.895 ;
        RECT 20.895 11.725 21.235 11.895 ;
        RECT 21.685 11.725 22.025 11.895 ;
        RECT 22.475 11.725 22.815 11.895 ;
        RECT 25.550 11.720 25.890 11.890 ;
        RECT 26.340 11.720 26.680 11.890 ;
        RECT 27.130 11.720 27.470 11.890 ;
        RECT 27.920 11.720 28.260 11.890 ;
        RECT 28.710 11.720 29.050 11.890 ;
        RECT 29.500 11.720 29.840 11.890 ;
        RECT 30.290 11.720 30.630 11.890 ;
        RECT 31.080 11.720 31.420 11.890 ;
        RECT 31.870 11.720 32.210 11.890 ;
        RECT 32.660 11.720 33.000 11.890 ;
        RECT 35.490 11.720 35.830 11.890 ;
        RECT 36.280 11.720 36.620 11.890 ;
        RECT 37.070 11.720 37.410 11.890 ;
        RECT 37.860 11.720 38.200 11.890 ;
        RECT 38.650 11.720 38.990 11.890 ;
        RECT 39.440 11.720 39.780 11.890 ;
        RECT 40.230 11.720 40.570 11.890 ;
        RECT 41.020 11.720 41.360 11.890 ;
        RECT 41.810 11.720 42.150 11.890 ;
        RECT 42.600 11.720 42.940 11.890 ;
        RECT 45.290 11.720 45.630 11.890 ;
        RECT 46.080 11.720 46.420 11.890 ;
        RECT 46.870 11.720 47.210 11.890 ;
        RECT 47.660 11.720 48.000 11.890 ;
        RECT 48.450 11.720 48.790 11.890 ;
        RECT 49.240 11.720 49.580 11.890 ;
        RECT 50.030 11.720 50.370 11.890 ;
        RECT 50.820 11.720 51.160 11.890 ;
        RECT 51.610 11.720 51.950 11.890 ;
        RECT 52.400 11.720 52.740 11.890 ;
        RECT 55.090 11.720 55.430 11.890 ;
        RECT 55.880 11.720 56.220 11.890 ;
        RECT 56.670 11.720 57.010 11.890 ;
        RECT 57.460 11.720 57.800 11.890 ;
        RECT 58.250 11.720 58.590 11.890 ;
        RECT 59.040 11.720 59.380 11.890 ;
        RECT 59.830 11.720 60.170 11.890 ;
        RECT 60.620 11.720 60.960 11.890 ;
        RECT 61.410 11.720 61.750 11.890 ;
        RECT 62.200 11.720 62.540 11.890 ;
        RECT 64.890 11.720 65.230 11.890 ;
        RECT 65.680 11.720 66.020 11.890 ;
        RECT 66.470 11.720 66.810 11.890 ;
        RECT 67.260 11.720 67.600 11.890 ;
        RECT 68.050 11.720 68.390 11.890 ;
        RECT 68.840 11.720 69.180 11.890 ;
        RECT 69.630 11.720 69.970 11.890 ;
        RECT 70.420 11.720 70.760 11.890 ;
        RECT 71.210 11.720 71.550 11.890 ;
        RECT 72.000 11.720 72.340 11.890 ;
        RECT 15.845 1.545 16.015 11.425 ;
        RECT 17.425 1.545 17.595 11.425 ;
        RECT 19.005 1.545 19.175 11.425 ;
        RECT 20.585 1.545 20.755 11.425 ;
        RECT 22.165 1.545 22.335 11.425 ;
        RECT 15.365 1.075 15.705 1.245 ;
        RECT 16.155 1.075 16.495 1.245 ;
        RECT 16.945 1.075 17.285 1.245 ;
        RECT 17.735 1.075 18.075 1.245 ;
        RECT 18.525 1.075 18.865 1.245 ;
        RECT 19.315 1.075 19.655 1.245 ;
        RECT 20.105 1.075 20.445 1.245 ;
        RECT 20.895 1.075 21.235 1.245 ;
        RECT 21.685 1.075 22.025 1.245 ;
        RECT 22.475 1.075 22.815 1.245 ;
        RECT 25.550 1.080 25.890 1.250 ;
        RECT 26.340 1.080 26.680 1.250 ;
        RECT 27.130 1.080 27.470 1.250 ;
        RECT 27.920 1.080 28.260 1.250 ;
        RECT 28.710 1.080 29.050 1.250 ;
        RECT 29.500 1.080 29.840 1.250 ;
        RECT 30.290 1.080 30.630 1.250 ;
        RECT 31.080 1.080 31.420 1.250 ;
        RECT 31.870 1.080 32.210 1.250 ;
        RECT 32.660 1.080 33.000 1.250 ;
        RECT 35.490 1.080 35.830 1.250 ;
        RECT 36.280 1.080 36.620 1.250 ;
        RECT 37.070 1.080 37.410 1.250 ;
        RECT 37.860 1.080 38.200 1.250 ;
        RECT 38.650 1.080 38.990 1.250 ;
        RECT 39.440 1.080 39.780 1.250 ;
        RECT 40.230 1.080 40.570 1.250 ;
        RECT 41.020 1.080 41.360 1.250 ;
        RECT 41.810 1.080 42.150 1.250 ;
        RECT 42.600 1.080 42.940 1.250 ;
        RECT 45.290 1.080 45.630 1.250 ;
        RECT 46.080 1.080 46.420 1.250 ;
        RECT 46.870 1.080 47.210 1.250 ;
        RECT 47.660 1.080 48.000 1.250 ;
        RECT 48.450 1.080 48.790 1.250 ;
        RECT 49.240 1.080 49.580 1.250 ;
        RECT 50.030 1.080 50.370 1.250 ;
        RECT 50.820 1.080 51.160 1.250 ;
        RECT 51.610 1.080 51.950 1.250 ;
        RECT 52.400 1.080 52.740 1.250 ;
        RECT 55.090 1.080 55.430 1.250 ;
        RECT 55.880 1.080 56.220 1.250 ;
        RECT 56.670 1.080 57.010 1.250 ;
        RECT 57.460 1.080 57.800 1.250 ;
        RECT 58.250 1.080 58.590 1.250 ;
        RECT 59.040 1.080 59.380 1.250 ;
        RECT 59.830 1.080 60.170 1.250 ;
        RECT 60.620 1.080 60.960 1.250 ;
        RECT 61.410 1.080 61.750 1.250 ;
        RECT 62.200 1.080 62.540 1.250 ;
        RECT 64.890 1.080 65.230 1.250 ;
        RECT 65.680 1.080 66.020 1.250 ;
        RECT 66.470 1.080 66.810 1.250 ;
        RECT 67.260 1.080 67.600 1.250 ;
        RECT 68.050 1.080 68.390 1.250 ;
        RECT 68.840 1.080 69.180 1.250 ;
        RECT 69.630 1.080 69.970 1.250 ;
        RECT 70.420 1.080 70.760 1.250 ;
        RECT 71.210 1.080 71.550 1.250 ;
        RECT 72.000 1.080 72.340 1.250 ;
      LAYER met1 ;
        RECT 15.305 140.555 15.765 140.785 ;
        RECT 16.095 140.555 16.555 140.785 ;
        RECT 16.885 140.555 17.345 140.785 ;
        RECT 17.675 140.555 18.135 140.785 ;
        RECT 18.465 140.555 18.925 140.785 ;
        RECT 19.255 140.555 19.715 140.785 ;
        RECT 20.045 140.555 20.505 140.785 ;
        RECT 20.835 140.555 21.295 140.785 ;
        RECT 21.625 140.555 22.085 140.785 ;
        RECT 22.415 140.555 22.875 140.785 ;
        RECT 25.490 140.550 25.950 140.780 ;
        RECT 26.280 140.550 26.740 140.780 ;
        RECT 27.070 140.550 27.530 140.780 ;
        RECT 27.860 140.550 28.320 140.780 ;
        RECT 28.650 140.550 29.110 140.780 ;
        RECT 29.440 140.550 29.900 140.780 ;
        RECT 30.230 140.550 30.690 140.780 ;
        RECT 31.020 140.550 31.480 140.780 ;
        RECT 31.810 140.550 32.270 140.780 ;
        RECT 32.600 140.550 33.060 140.780 ;
        RECT 35.430 140.550 35.890 140.780 ;
        RECT 36.220 140.550 36.680 140.780 ;
        RECT 37.010 140.550 37.470 140.780 ;
        RECT 37.800 140.550 38.260 140.780 ;
        RECT 38.590 140.550 39.050 140.780 ;
        RECT 39.380 140.550 39.840 140.780 ;
        RECT 40.170 140.550 40.630 140.780 ;
        RECT 40.960 140.550 41.420 140.780 ;
        RECT 41.750 140.550 42.210 140.780 ;
        RECT 42.540 140.550 43.000 140.780 ;
        RECT 45.230 140.550 45.690 140.780 ;
        RECT 46.020 140.550 46.480 140.780 ;
        RECT 46.810 140.550 47.270 140.780 ;
        RECT 47.600 140.550 48.060 140.780 ;
        RECT 48.390 140.550 48.850 140.780 ;
        RECT 49.180 140.550 49.640 140.780 ;
        RECT 49.970 140.550 50.430 140.780 ;
        RECT 50.760 140.550 51.220 140.780 ;
        RECT 51.550 140.550 52.010 140.780 ;
        RECT 52.340 140.550 52.800 140.780 ;
        RECT 55.030 140.550 55.490 140.780 ;
        RECT 55.820 140.550 56.280 140.780 ;
        RECT 56.610 140.550 57.070 140.780 ;
        RECT 57.400 140.550 57.860 140.780 ;
        RECT 58.190 140.550 58.650 140.780 ;
        RECT 58.980 140.550 59.440 140.780 ;
        RECT 59.770 140.550 60.230 140.780 ;
        RECT 60.560 140.550 61.020 140.780 ;
        RECT 61.350 140.550 61.810 140.780 ;
        RECT 62.140 140.550 62.600 140.780 ;
        RECT 64.830 140.550 65.290 140.780 ;
        RECT 65.620 140.550 66.080 140.780 ;
        RECT 66.410 140.550 66.870 140.780 ;
        RECT 67.200 140.550 67.660 140.780 ;
        RECT 67.990 140.550 68.450 140.780 ;
        RECT 68.780 140.550 69.240 140.780 ;
        RECT 69.570 140.550 70.030 140.780 ;
        RECT 70.360 140.550 70.820 140.780 ;
        RECT 71.150 140.550 71.610 140.780 ;
        RECT 71.940 140.550 72.400 140.780 ;
        RECT 15.815 131.360 16.045 140.345 ;
        RECT 17.395 131.360 17.625 140.345 ;
        RECT 18.975 131.360 19.215 140.345 ;
        RECT 15.720 130.710 16.120 131.360 ;
        RECT 17.310 130.710 17.710 131.360 ;
        RECT 18.890 130.710 19.290 131.360 ;
        RECT 20.555 131.350 20.785 140.345 ;
        RECT 22.135 131.350 22.365 140.345 ;
        RECT 15.815 130.345 16.045 130.710 ;
        RECT 17.395 130.345 17.625 130.710 ;
        RECT 18.975 130.345 19.215 130.710 ;
        RECT 20.450 130.700 20.850 131.350 ;
        RECT 22.030 130.700 22.430 131.350 ;
        RECT 20.555 130.345 20.785 130.700 ;
        RECT 22.135 130.345 22.365 130.700 ;
        RECT 13.980 129.360 22.900 130.160 ;
        RECT 25.490 130.125 25.950 130.140 ;
        RECT 26.280 130.130 26.740 130.140 ;
        RECT 27.070 130.130 27.530 130.140 ;
        RECT 27.860 130.130 28.320 130.140 ;
        RECT 28.650 130.130 29.110 130.140 ;
        RECT 29.440 130.130 29.900 130.140 ;
        RECT 30.230 130.130 30.690 130.140 ;
        RECT 31.020 130.130 31.480 130.140 ;
        RECT 31.810 130.130 32.270 130.140 ;
        RECT 32.600 130.130 33.060 130.140 ;
        RECT 35.430 130.130 35.890 130.140 ;
        RECT 36.220 130.130 36.680 130.140 ;
        RECT 37.010 130.130 37.470 130.140 ;
        RECT 37.800 130.130 38.260 130.140 ;
        RECT 38.590 130.130 39.050 130.140 ;
        RECT 39.380 130.130 39.840 130.140 ;
        RECT 40.170 130.130 40.630 130.140 ;
        RECT 40.960 130.130 41.420 130.140 ;
        RECT 41.750 130.130 42.210 130.140 ;
        RECT 42.540 130.130 43.000 130.140 ;
        RECT 45.230 130.130 45.690 130.140 ;
        RECT 46.020 130.130 46.480 130.140 ;
        RECT 46.810 130.130 47.270 130.140 ;
        RECT 47.600 130.130 48.060 130.140 ;
        RECT 48.390 130.130 48.850 130.140 ;
        RECT 49.180 130.130 49.640 130.140 ;
        RECT 49.970 130.130 50.430 130.140 ;
        RECT 50.760 130.130 51.220 130.140 ;
        RECT 51.550 130.130 52.010 130.140 ;
        RECT 52.340 130.130 52.800 130.140 ;
        RECT 55.030 130.130 55.490 130.140 ;
        RECT 55.820 130.130 56.280 130.140 ;
        RECT 56.610 130.130 57.070 130.140 ;
        RECT 57.400 130.130 57.860 130.140 ;
        RECT 58.190 130.130 58.650 130.140 ;
        RECT 58.980 130.130 59.440 130.140 ;
        RECT 59.770 130.130 60.230 130.140 ;
        RECT 60.560 130.130 61.020 130.140 ;
        RECT 61.350 130.130 61.810 130.140 ;
        RECT 62.140 130.130 62.600 130.140 ;
        RECT 64.830 130.130 65.290 130.140 ;
        RECT 65.620 130.130 66.080 130.140 ;
        RECT 66.410 130.130 66.870 130.140 ;
        RECT 67.200 130.130 67.660 130.140 ;
        RECT 67.990 130.130 68.450 130.140 ;
        RECT 68.780 130.130 69.240 130.140 ;
        RECT 69.570 130.130 70.030 130.140 ;
        RECT 70.360 130.130 70.820 130.140 ;
        RECT 71.150 130.130 71.610 130.140 ;
        RECT 71.940 130.130 72.400 130.140 ;
        RECT 26.215 130.125 72.400 130.130 ;
        RECT 23.875 130.080 72.400 130.125 ;
        RECT 23.860 129.360 72.400 130.080 ;
        RECT 13.980 103.630 14.780 129.360 ;
        RECT 23.860 129.355 26.215 129.360 ;
        RECT 15.815 128.670 16.045 129.165 ;
        RECT 17.395 128.680 17.625 129.165 ;
        RECT 18.975 128.680 19.205 129.165 ;
        RECT 20.555 128.690 20.785 129.165 ;
        RECT 22.135 128.690 22.365 129.165 ;
        RECT 15.730 128.020 16.130 128.670 ;
        RECT 17.310 128.030 17.710 128.680 ;
        RECT 18.880 128.030 19.280 128.680 ;
        RECT 20.460 128.040 20.860 128.690 ;
        RECT 22.030 128.040 22.430 128.690 ;
        RECT 23.860 128.470 24.660 129.355 ;
        RECT 15.815 119.165 16.045 128.020 ;
        RECT 17.395 119.165 17.625 128.030 ;
        RECT 18.975 119.165 19.205 128.030 ;
        RECT 20.555 119.165 20.785 128.040 ;
        RECT 22.135 119.165 22.365 128.040 ;
        RECT 15.305 118.725 15.765 118.955 ;
        RECT 16.095 118.725 16.555 118.955 ;
        RECT 16.885 118.725 17.345 118.955 ;
        RECT 17.675 118.725 18.135 118.955 ;
        RECT 18.465 118.725 18.925 118.955 ;
        RECT 19.255 118.725 19.715 118.955 ;
        RECT 20.045 118.725 20.505 118.955 ;
        RECT 20.835 118.725 21.295 118.955 ;
        RECT 21.625 118.725 22.085 118.955 ;
        RECT 22.415 118.725 22.875 118.955 ;
        RECT 16.560 116.790 17.020 117.020 ;
        RECT 17.350 116.790 17.810 117.020 ;
        RECT 20.045 116.795 20.505 117.025 ;
        RECT 20.835 116.795 21.295 117.025 ;
        RECT 21.625 116.795 22.085 117.025 ;
        RECT 22.415 116.795 22.875 117.025 ;
        RECT 17.070 113.580 17.300 116.580 ;
        RECT 16.980 112.930 17.380 113.580 ;
        RECT 17.070 112.580 17.300 112.930 ;
        RECT 13.960 102.610 14.780 103.630 ;
        RECT 13.980 94.870 14.780 102.610 ;
        RECT 15.430 112.120 17.880 112.380 ;
        RECT 15.430 110.530 15.690 112.120 ;
        RECT 15.430 110.270 18.080 110.530 ;
        RECT 15.430 103.390 15.690 110.270 ;
        RECT 16.240 110.020 16.500 110.270 ;
        RECT 17.820 110.020 18.080 110.270 ;
        RECT 16.240 109.860 16.505 110.020 ;
        RECT 16.170 109.210 16.570 109.860 ;
        RECT 17.820 109.850 18.085 110.020 ;
        RECT 16.275 109.020 16.505 109.210 ;
        RECT 17.760 109.200 18.160 109.850 ;
        RECT 17.855 109.020 18.085 109.200 ;
        RECT 16.555 108.580 17.805 108.810 ;
        RECT 16.850 106.930 17.390 108.580 ;
        RECT 20.555 107.620 20.785 116.585 ;
        RECT 22.135 107.630 22.365 116.585 ;
        RECT 23.875 107.770 24.645 128.470 ;
        RECT 25.490 118.730 25.950 118.960 ;
        RECT 26.280 118.730 26.740 118.960 ;
        RECT 27.070 118.730 27.530 118.960 ;
        RECT 27.860 118.730 28.320 118.960 ;
        RECT 28.650 118.730 29.110 118.960 ;
        RECT 29.440 118.730 29.900 118.960 ;
        RECT 30.230 118.730 30.690 118.960 ;
        RECT 31.020 118.730 31.480 118.960 ;
        RECT 31.810 118.730 32.270 118.960 ;
        RECT 32.600 118.730 33.060 118.960 ;
        RECT 35.430 118.730 35.890 118.960 ;
        RECT 36.220 118.730 36.680 118.960 ;
        RECT 37.010 118.730 37.470 118.960 ;
        RECT 37.800 118.730 38.260 118.960 ;
        RECT 38.590 118.730 39.050 118.960 ;
        RECT 39.380 118.730 39.840 118.960 ;
        RECT 40.170 118.730 40.630 118.960 ;
        RECT 40.960 118.730 41.420 118.960 ;
        RECT 41.750 118.730 42.210 118.960 ;
        RECT 42.540 118.730 43.000 118.960 ;
        RECT 45.230 118.730 45.690 118.960 ;
        RECT 46.020 118.730 46.480 118.960 ;
        RECT 46.810 118.730 47.270 118.960 ;
        RECT 47.600 118.730 48.060 118.960 ;
        RECT 48.390 118.730 48.850 118.960 ;
        RECT 49.180 118.730 49.640 118.960 ;
        RECT 49.970 118.730 50.430 118.960 ;
        RECT 50.760 118.730 51.220 118.960 ;
        RECT 51.550 118.730 52.010 118.960 ;
        RECT 52.340 118.730 52.800 118.960 ;
        RECT 55.030 118.730 55.490 118.960 ;
        RECT 55.820 118.730 56.280 118.960 ;
        RECT 56.610 118.730 57.070 118.960 ;
        RECT 57.400 118.730 57.860 118.960 ;
        RECT 58.190 118.730 58.650 118.960 ;
        RECT 58.980 118.730 59.440 118.960 ;
        RECT 59.770 118.730 60.230 118.960 ;
        RECT 60.560 118.730 61.020 118.960 ;
        RECT 61.350 118.730 61.810 118.960 ;
        RECT 62.140 118.730 62.600 118.960 ;
        RECT 64.830 118.730 65.290 118.960 ;
        RECT 65.620 118.730 66.080 118.960 ;
        RECT 66.410 118.730 66.870 118.960 ;
        RECT 67.200 118.730 67.660 118.960 ;
        RECT 67.990 118.730 68.450 118.960 ;
        RECT 68.780 118.730 69.240 118.960 ;
        RECT 69.570 118.730 70.030 118.960 ;
        RECT 70.360 118.730 70.820 118.960 ;
        RECT 71.150 118.730 71.610 118.960 ;
        RECT 71.940 118.730 72.400 118.960 ;
        RECT 25.490 118.190 25.950 118.420 ;
        RECT 26.280 118.190 26.740 118.420 ;
        RECT 27.070 118.190 27.530 118.420 ;
        RECT 27.860 118.190 28.320 118.420 ;
        RECT 28.650 118.190 29.110 118.420 ;
        RECT 29.440 118.190 29.900 118.420 ;
        RECT 30.230 118.190 30.690 118.420 ;
        RECT 31.020 118.190 31.480 118.420 ;
        RECT 31.810 118.190 32.270 118.420 ;
        RECT 32.600 118.190 33.060 118.420 ;
        RECT 35.430 118.190 35.890 118.420 ;
        RECT 36.220 118.190 36.680 118.420 ;
        RECT 37.010 118.190 37.470 118.420 ;
        RECT 37.800 118.190 38.260 118.420 ;
        RECT 38.590 118.190 39.050 118.420 ;
        RECT 39.380 118.190 39.840 118.420 ;
        RECT 40.170 118.190 40.630 118.420 ;
        RECT 40.960 118.190 41.420 118.420 ;
        RECT 41.750 118.190 42.210 118.420 ;
        RECT 42.540 118.190 43.000 118.420 ;
        RECT 45.230 118.190 45.690 118.420 ;
        RECT 46.020 118.190 46.480 118.420 ;
        RECT 46.810 118.190 47.270 118.420 ;
        RECT 47.600 118.190 48.060 118.420 ;
        RECT 48.390 118.190 48.850 118.420 ;
        RECT 49.180 118.190 49.640 118.420 ;
        RECT 49.970 118.190 50.430 118.420 ;
        RECT 50.760 118.190 51.220 118.420 ;
        RECT 51.550 118.190 52.010 118.420 ;
        RECT 52.340 118.190 52.800 118.420 ;
        RECT 55.030 118.190 55.490 118.420 ;
        RECT 55.820 118.190 56.280 118.420 ;
        RECT 56.610 118.190 57.070 118.420 ;
        RECT 57.400 118.190 57.860 118.420 ;
        RECT 58.190 118.190 58.650 118.420 ;
        RECT 58.980 118.190 59.440 118.420 ;
        RECT 59.770 118.190 60.230 118.420 ;
        RECT 60.560 118.190 61.020 118.420 ;
        RECT 61.350 118.190 61.810 118.420 ;
        RECT 62.140 118.190 62.600 118.420 ;
        RECT 64.830 118.190 65.290 118.420 ;
        RECT 65.620 118.190 66.080 118.420 ;
        RECT 66.410 118.190 66.870 118.420 ;
        RECT 67.200 118.190 67.660 118.420 ;
        RECT 67.990 118.190 68.450 118.420 ;
        RECT 68.780 118.190 69.240 118.420 ;
        RECT 69.570 118.190 70.030 118.420 ;
        RECT 70.360 118.190 70.820 118.420 ;
        RECT 71.150 118.190 71.610 118.420 ;
        RECT 71.940 118.190 72.400 118.420 ;
        RECT 25.490 107.770 25.950 107.780 ;
        RECT 26.280 107.770 26.740 107.780 ;
        RECT 27.070 107.770 27.530 107.780 ;
        RECT 27.860 107.770 28.320 107.780 ;
        RECT 28.650 107.770 29.110 107.780 ;
        RECT 29.440 107.770 29.900 107.780 ;
        RECT 30.230 107.770 30.690 107.780 ;
        RECT 31.020 107.770 31.480 107.780 ;
        RECT 31.810 107.770 32.270 107.780 ;
        RECT 32.600 107.770 33.060 107.780 ;
        RECT 35.430 107.770 35.890 107.780 ;
        RECT 36.220 107.770 36.680 107.780 ;
        RECT 37.010 107.770 37.470 107.780 ;
        RECT 37.800 107.770 38.260 107.780 ;
        RECT 38.590 107.770 39.050 107.780 ;
        RECT 39.380 107.770 39.840 107.780 ;
        RECT 40.170 107.770 40.630 107.780 ;
        RECT 40.960 107.770 41.420 107.780 ;
        RECT 41.750 107.770 42.210 107.780 ;
        RECT 42.540 107.770 43.000 107.780 ;
        RECT 45.230 107.770 45.690 107.780 ;
        RECT 46.020 107.770 46.480 107.780 ;
        RECT 46.810 107.770 47.270 107.780 ;
        RECT 47.600 107.770 48.060 107.780 ;
        RECT 48.390 107.770 48.850 107.780 ;
        RECT 49.180 107.770 49.640 107.780 ;
        RECT 49.970 107.770 50.430 107.780 ;
        RECT 50.760 107.770 51.220 107.780 ;
        RECT 51.550 107.770 52.010 107.780 ;
        RECT 52.340 107.770 52.800 107.780 ;
        RECT 55.030 107.770 55.490 107.780 ;
        RECT 55.820 107.770 56.280 107.780 ;
        RECT 56.610 107.770 57.070 107.780 ;
        RECT 57.400 107.770 57.860 107.780 ;
        RECT 58.190 107.770 58.650 107.780 ;
        RECT 58.980 107.770 59.440 107.780 ;
        RECT 59.770 107.770 60.230 107.780 ;
        RECT 60.560 107.770 61.020 107.780 ;
        RECT 61.350 107.770 61.810 107.780 ;
        RECT 62.140 107.770 62.600 107.780 ;
        RECT 64.830 107.770 65.290 107.780 ;
        RECT 65.620 107.770 66.080 107.780 ;
        RECT 66.410 107.770 66.870 107.780 ;
        RECT 67.200 107.770 67.660 107.780 ;
        RECT 67.990 107.770 68.450 107.780 ;
        RECT 68.780 107.770 69.240 107.780 ;
        RECT 69.570 107.770 70.030 107.780 ;
        RECT 70.360 107.770 70.820 107.780 ;
        RECT 71.150 107.770 71.610 107.780 ;
        RECT 71.940 107.770 72.400 107.780 ;
        RECT 20.470 106.970 20.870 107.620 ;
        RECT 22.070 106.980 22.470 107.630 ;
        RECT 23.875 107.000 72.400 107.770 ;
        RECT 16.820 106.390 17.420 106.930 ;
        RECT 20.555 106.585 20.785 106.970 ;
        RECT 22.135 106.585 22.365 106.980 ;
        RECT 16.850 103.910 17.390 106.390 ;
        RECT 20.030 106.120 22.900 106.400 ;
        RECT 20.410 105.510 20.860 106.120 ;
        RECT 20.210 104.900 20.860 105.510 ;
        RECT 16.580 103.390 16.810 103.760 ;
        RECT 15.430 103.130 16.810 103.390 ;
        RECT 15.430 100.680 15.690 103.130 ;
        RECT 16.580 102.760 16.810 103.130 ;
        RECT 16.860 102.370 17.320 102.600 ;
        RECT 20.410 102.535 20.860 104.900 ;
        RECT 18.195 102.085 20.860 102.535 ;
        RECT 15.430 100.660 17.310 100.680 ;
        RECT 15.430 100.430 17.320 100.660 ;
        RECT 15.430 100.420 17.310 100.430 ;
        RECT 17.370 98.945 17.600 100.270 ;
        RECT 18.195 98.945 18.645 102.085 ;
        RECT 20.410 101.690 20.860 102.085 ;
        RECT 19.520 101.410 22.390 101.690 ;
        RECT 20.065 100.740 20.295 101.270 ;
        RECT 21.645 100.740 21.875 101.270 ;
        RECT 19.970 100.090 20.370 100.740 ;
        RECT 21.560 100.090 21.960 100.740 ;
        RECT 17.370 98.495 18.645 98.945 ;
        RECT 17.370 96.270 17.600 98.495 ;
        RECT 20.065 96.270 20.295 100.090 ;
        RECT 21.645 96.270 21.875 100.090 ;
        RECT 16.860 95.880 17.320 96.110 ;
        RECT 19.555 95.880 20.015 96.110 ;
        RECT 20.345 95.880 20.805 96.110 ;
        RECT 21.135 95.880 21.595 96.110 ;
        RECT 21.925 95.880 22.385 96.110 ;
        RECT 13.595 94.200 22.870 94.870 ;
        RECT 13.595 93.920 22.880 94.200 ;
        RECT 3.615 80.660 4.075 80.890 ;
        RECT 4.405 80.660 4.865 80.890 ;
        RECT 5.195 80.660 5.655 80.890 ;
        RECT 5.985 80.660 6.445 80.890 ;
        RECT 6.775 80.660 7.235 80.890 ;
        RECT 8.905 80.660 9.365 80.890 ;
        RECT 9.695 80.660 10.155 80.890 ;
        RECT 10.485 80.660 10.945 80.890 ;
        RECT 11.275 80.660 11.735 80.890 ;
        RECT 12.065 80.660 12.525 80.890 ;
        RECT 4.125 79.055 4.355 80.450 ;
        RECT 5.705 79.055 5.935 80.450 ;
        RECT 7.285 79.055 7.515 80.450 ;
        RECT 8.625 79.055 8.855 80.450 ;
        RECT 10.205 79.055 10.435 80.450 ;
        RECT 11.785 79.055 12.015 80.450 ;
        RECT 4.045 78.455 4.435 79.055 ;
        RECT 5.625 78.455 6.015 79.055 ;
        RECT 7.205 78.455 7.595 79.055 ;
        RECT 8.545 78.825 8.935 79.055 ;
        RECT 4.125 78.450 4.355 78.455 ;
        RECT 5.705 78.450 5.935 78.455 ;
        RECT 7.285 78.450 7.515 78.455 ;
        RECT 8.015 78.445 8.935 78.825 ;
        RECT 10.125 78.455 10.515 79.055 ;
        RECT 11.705 78.455 12.095 79.055 ;
        RECT 13.595 78.635 14.545 93.920 ;
        RECT 15.815 93.240 16.045 93.760 ;
        RECT 17.395 93.240 17.625 93.760 ;
        RECT 15.730 92.590 16.130 93.240 ;
        RECT 17.300 92.590 17.700 93.240 ;
        RECT 18.975 93.230 19.205 93.760 ;
        RECT 20.555 93.230 20.785 93.760 ;
        RECT 15.815 83.760 16.045 92.590 ;
        RECT 17.395 83.760 17.625 92.590 ;
        RECT 18.880 92.580 19.280 93.230 ;
        RECT 20.470 92.580 20.870 93.230 ;
        RECT 22.135 93.220 22.365 93.760 ;
        RECT 18.975 83.760 19.205 92.580 ;
        RECT 20.555 83.760 20.785 92.580 ;
        RECT 22.060 92.570 22.460 93.220 ;
        RECT 22.135 83.760 22.365 92.570 ;
        RECT 23.875 83.610 24.645 107.000 ;
        RECT 25.490 96.370 25.950 96.600 ;
        RECT 26.280 96.370 26.740 96.600 ;
        RECT 27.070 96.370 27.530 96.600 ;
        RECT 27.860 96.370 28.320 96.600 ;
        RECT 28.650 96.370 29.110 96.600 ;
        RECT 29.440 96.370 29.900 96.600 ;
        RECT 30.230 96.370 30.690 96.600 ;
        RECT 31.020 96.370 31.480 96.600 ;
        RECT 31.810 96.370 32.270 96.600 ;
        RECT 32.600 96.370 33.060 96.600 ;
        RECT 35.430 96.370 35.890 96.600 ;
        RECT 36.220 96.370 36.680 96.600 ;
        RECT 37.010 96.370 37.470 96.600 ;
        RECT 37.800 96.370 38.260 96.600 ;
        RECT 38.590 96.370 39.050 96.600 ;
        RECT 39.380 96.370 39.840 96.600 ;
        RECT 40.170 96.370 40.630 96.600 ;
        RECT 40.960 96.370 41.420 96.600 ;
        RECT 41.750 96.370 42.210 96.600 ;
        RECT 42.540 96.370 43.000 96.600 ;
        RECT 45.230 96.370 45.690 96.600 ;
        RECT 46.020 96.370 46.480 96.600 ;
        RECT 46.810 96.370 47.270 96.600 ;
        RECT 47.600 96.370 48.060 96.600 ;
        RECT 48.390 96.370 48.850 96.600 ;
        RECT 49.180 96.370 49.640 96.600 ;
        RECT 49.970 96.370 50.430 96.600 ;
        RECT 50.760 96.370 51.220 96.600 ;
        RECT 51.550 96.370 52.010 96.600 ;
        RECT 52.340 96.370 52.800 96.600 ;
        RECT 55.030 96.370 55.490 96.600 ;
        RECT 55.820 96.370 56.280 96.600 ;
        RECT 56.610 96.370 57.070 96.600 ;
        RECT 57.400 96.370 57.860 96.600 ;
        RECT 58.190 96.370 58.650 96.600 ;
        RECT 58.980 96.370 59.440 96.600 ;
        RECT 59.770 96.370 60.230 96.600 ;
        RECT 60.560 96.370 61.020 96.600 ;
        RECT 61.350 96.370 61.810 96.600 ;
        RECT 62.140 96.370 62.600 96.600 ;
        RECT 64.830 96.370 65.290 96.600 ;
        RECT 65.620 96.370 66.080 96.600 ;
        RECT 66.410 96.370 66.870 96.600 ;
        RECT 67.200 96.370 67.660 96.600 ;
        RECT 67.990 96.370 68.450 96.600 ;
        RECT 68.780 96.370 69.240 96.600 ;
        RECT 69.570 96.370 70.030 96.600 ;
        RECT 70.360 96.370 70.820 96.600 ;
        RECT 71.150 96.370 71.610 96.600 ;
        RECT 71.940 96.370 72.400 96.600 ;
        RECT 25.495 93.935 25.955 94.165 ;
        RECT 26.285 93.935 26.745 94.165 ;
        RECT 27.075 93.935 27.535 94.165 ;
        RECT 27.865 93.935 28.325 94.165 ;
        RECT 28.655 93.935 29.115 94.165 ;
        RECT 29.445 93.935 29.905 94.165 ;
        RECT 30.235 93.935 30.695 94.165 ;
        RECT 31.025 93.935 31.485 94.165 ;
        RECT 31.815 93.935 32.275 94.165 ;
        RECT 32.605 93.935 33.065 94.165 ;
        RECT 35.435 93.935 35.895 94.165 ;
        RECT 36.225 93.935 36.685 94.165 ;
        RECT 37.015 93.935 37.475 94.165 ;
        RECT 37.805 93.935 38.265 94.165 ;
        RECT 38.595 93.935 39.055 94.165 ;
        RECT 39.385 93.935 39.845 94.165 ;
        RECT 40.175 93.935 40.635 94.165 ;
        RECT 40.965 93.935 41.425 94.165 ;
        RECT 41.755 93.935 42.215 94.165 ;
        RECT 42.545 93.935 43.005 94.165 ;
        RECT 45.235 93.935 45.695 94.165 ;
        RECT 46.025 93.935 46.485 94.165 ;
        RECT 46.815 93.935 47.275 94.165 ;
        RECT 47.605 93.935 48.065 94.165 ;
        RECT 48.395 93.935 48.855 94.165 ;
        RECT 49.185 93.935 49.645 94.165 ;
        RECT 49.975 93.935 50.435 94.165 ;
        RECT 50.765 93.935 51.225 94.165 ;
        RECT 51.555 93.935 52.015 94.165 ;
        RECT 52.345 93.935 52.805 94.165 ;
        RECT 55.035 93.935 55.495 94.165 ;
        RECT 55.825 93.935 56.285 94.165 ;
        RECT 56.615 93.935 57.075 94.165 ;
        RECT 57.405 93.935 57.865 94.165 ;
        RECT 58.195 93.935 58.655 94.165 ;
        RECT 58.985 93.935 59.445 94.165 ;
        RECT 59.775 93.935 60.235 94.165 ;
        RECT 60.565 93.935 61.025 94.165 ;
        RECT 61.355 93.935 61.815 94.165 ;
        RECT 62.145 93.935 62.605 94.165 ;
        RECT 64.835 93.935 65.295 94.165 ;
        RECT 65.625 93.935 66.085 94.165 ;
        RECT 66.415 93.935 66.875 94.165 ;
        RECT 67.205 93.935 67.665 94.165 ;
        RECT 67.995 93.935 68.455 94.165 ;
        RECT 68.785 93.935 69.245 94.165 ;
        RECT 69.575 93.935 70.035 94.165 ;
        RECT 70.365 93.935 70.825 94.165 ;
        RECT 71.155 93.935 71.615 94.165 ;
        RECT 71.945 93.935 72.405 94.165 ;
        RECT 25.495 83.610 25.955 83.615 ;
        RECT 26.285 83.610 26.745 83.615 ;
        RECT 27.075 83.610 27.535 83.615 ;
        RECT 27.865 83.610 28.325 83.615 ;
        RECT 28.655 83.610 29.115 83.615 ;
        RECT 29.445 83.610 29.905 83.615 ;
        RECT 30.235 83.610 30.695 83.615 ;
        RECT 31.025 83.610 31.485 83.615 ;
        RECT 31.815 83.610 32.275 83.615 ;
        RECT 32.605 83.610 33.065 83.615 ;
        RECT 35.435 83.610 35.895 83.615 ;
        RECT 36.225 83.610 36.685 83.615 ;
        RECT 37.015 83.610 37.475 83.615 ;
        RECT 37.805 83.610 38.265 83.615 ;
        RECT 38.595 83.610 39.055 83.615 ;
        RECT 39.385 83.610 39.845 83.615 ;
        RECT 40.175 83.610 40.635 83.615 ;
        RECT 40.965 83.610 41.425 83.615 ;
        RECT 41.755 83.610 42.215 83.615 ;
        RECT 42.545 83.610 43.005 83.615 ;
        RECT 45.235 83.610 45.695 83.615 ;
        RECT 46.025 83.610 46.485 83.615 ;
        RECT 46.815 83.610 47.275 83.615 ;
        RECT 47.605 83.610 48.065 83.615 ;
        RECT 48.395 83.610 48.855 83.615 ;
        RECT 49.185 83.610 49.645 83.615 ;
        RECT 49.975 83.610 50.435 83.615 ;
        RECT 50.765 83.610 51.225 83.615 ;
        RECT 51.555 83.610 52.015 83.615 ;
        RECT 52.345 83.610 52.805 83.615 ;
        RECT 55.035 83.610 55.495 83.615 ;
        RECT 55.825 83.610 56.285 83.615 ;
        RECT 56.615 83.610 57.075 83.615 ;
        RECT 57.405 83.610 57.865 83.615 ;
        RECT 58.195 83.610 58.655 83.615 ;
        RECT 58.985 83.610 59.445 83.615 ;
        RECT 59.775 83.610 60.235 83.615 ;
        RECT 60.565 83.610 61.025 83.615 ;
        RECT 61.355 83.610 61.815 83.615 ;
        RECT 62.145 83.610 62.605 83.615 ;
        RECT 64.835 83.610 65.295 83.615 ;
        RECT 65.625 83.610 66.085 83.615 ;
        RECT 66.415 83.610 66.875 83.615 ;
        RECT 67.205 83.610 67.665 83.615 ;
        RECT 67.995 83.610 68.455 83.615 ;
        RECT 68.785 83.610 69.245 83.615 ;
        RECT 69.575 83.610 70.035 83.615 ;
        RECT 70.365 83.610 70.825 83.615 ;
        RECT 71.155 83.610 71.615 83.615 ;
        RECT 71.945 83.610 72.405 83.615 ;
        RECT 15.305 83.370 15.765 83.600 ;
        RECT 16.095 83.370 16.555 83.600 ;
        RECT 16.885 83.370 17.345 83.600 ;
        RECT 17.675 83.370 18.135 83.600 ;
        RECT 18.465 83.370 18.925 83.600 ;
        RECT 19.255 83.370 19.715 83.600 ;
        RECT 20.045 83.370 20.505 83.600 ;
        RECT 20.835 83.370 21.295 83.600 ;
        RECT 21.625 83.370 22.085 83.600 ;
        RECT 22.415 83.370 22.875 83.600 ;
        RECT 23.875 83.385 72.405 83.610 ;
        RECT 23.875 83.085 72.400 83.385 ;
        RECT 23.875 82.855 72.405 83.085 ;
        RECT 23.875 82.840 72.400 82.855 ;
        RECT 17.985 80.080 18.445 80.310 ;
        RECT 18.775 80.080 19.235 80.310 ;
        RECT 21.065 80.080 21.525 80.310 ;
        RECT 21.855 80.080 22.315 80.310 ;
        RECT 10.205 78.450 10.435 78.455 ;
        RECT 11.785 78.450 12.015 78.455 ;
        RECT 8.015 78.255 8.375 78.445 ;
        RECT 3.615 78.015 8.375 78.255 ;
        RECT 8.905 78.015 12.525 78.255 ;
        RECT 3.615 78.010 4.075 78.015 ;
        RECT 4.405 78.010 4.865 78.015 ;
        RECT 5.195 78.010 5.655 78.015 ;
        RECT 5.985 78.010 6.445 78.015 ;
        RECT 6.775 78.010 7.235 78.015 ;
        RECT 8.905 78.010 9.365 78.015 ;
        RECT 9.695 78.010 10.155 78.015 ;
        RECT 10.485 78.010 10.945 78.015 ;
        RECT 11.275 78.010 11.735 78.015 ;
        RECT 12.065 78.010 12.525 78.015 ;
        RECT 8.905 77.605 9.265 78.010 ;
        RECT 13.595 77.685 17.035 78.635 ;
        RECT 0.985 74.775 1.215 75.315 ;
        RECT 0.895 73.615 1.305 74.775 ;
        RECT 0.985 65.315 1.215 73.615 ;
        RECT 2.175 65.705 2.405 75.315 ;
        RECT 3.365 74.775 3.595 75.315 ;
        RECT 3.285 73.615 3.695 74.775 ;
        RECT 2.115 65.315 2.475 65.705 ;
        RECT 3.365 65.315 3.595 73.615 ;
        RECT 4.555 65.705 4.785 75.315 ;
        RECT 5.745 74.775 5.975 75.315 ;
        RECT 5.665 73.615 6.075 74.775 ;
        RECT 4.495 65.315 4.855 65.705 ;
        RECT 5.745 65.315 5.975 73.615 ;
        RECT 6.935 65.705 7.165 75.315 ;
        RECT 8.835 65.705 9.065 75.315 ;
        RECT 10.025 74.775 10.255 75.315 ;
        RECT 9.945 73.615 10.355 74.775 ;
        RECT 6.875 65.315 7.235 65.705 ;
        RECT 8.775 65.315 9.135 65.705 ;
        RECT 10.025 65.315 10.255 73.615 ;
        RECT 11.215 65.705 11.445 75.315 ;
        RECT 12.405 74.775 12.635 75.315 ;
        RECT 12.325 73.615 12.735 74.775 ;
        RECT 11.155 65.315 11.515 65.705 ;
        RECT 12.405 65.315 12.635 73.615 ;
        RECT 13.595 65.705 13.825 75.315 ;
        RECT 14.785 74.775 15.015 75.315 ;
        RECT 14.705 73.615 15.115 74.775 ;
        RECT 13.535 65.315 13.895 65.705 ;
        RECT 14.785 65.315 15.015 73.615 ;
        RECT 16.085 68.865 17.035 77.685 ;
        RECT 18.495 70.470 18.725 79.870 ;
        RECT 21.575 70.470 21.805 79.870 ;
        RECT 25.495 72.305 25.955 72.535 ;
        RECT 26.285 72.305 26.745 72.535 ;
        RECT 27.075 72.305 27.535 72.535 ;
        RECT 27.865 72.305 28.325 72.535 ;
        RECT 28.655 72.305 29.115 72.535 ;
        RECT 29.445 72.305 29.905 72.535 ;
        RECT 30.235 72.305 30.695 72.535 ;
        RECT 31.025 72.305 31.485 72.535 ;
        RECT 31.815 72.305 32.275 72.535 ;
        RECT 32.605 72.305 33.065 72.535 ;
        RECT 35.435 72.305 35.895 72.535 ;
        RECT 36.225 72.305 36.685 72.535 ;
        RECT 37.015 72.305 37.475 72.535 ;
        RECT 37.805 72.305 38.265 72.535 ;
        RECT 38.595 72.305 39.055 72.535 ;
        RECT 39.385 72.305 39.845 72.535 ;
        RECT 40.175 72.305 40.635 72.535 ;
        RECT 40.965 72.305 41.425 72.535 ;
        RECT 41.755 72.305 42.215 72.535 ;
        RECT 42.545 72.305 43.005 72.535 ;
        RECT 45.235 72.305 45.695 72.535 ;
        RECT 46.025 72.305 46.485 72.535 ;
        RECT 46.815 72.305 47.275 72.535 ;
        RECT 47.605 72.305 48.065 72.535 ;
        RECT 48.395 72.305 48.855 72.535 ;
        RECT 49.185 72.305 49.645 72.535 ;
        RECT 49.975 72.305 50.435 72.535 ;
        RECT 50.765 72.305 51.225 72.535 ;
        RECT 51.555 72.305 52.015 72.535 ;
        RECT 52.345 72.305 52.805 72.535 ;
        RECT 55.035 72.305 55.495 72.535 ;
        RECT 55.825 72.305 56.285 72.535 ;
        RECT 56.615 72.305 57.075 72.535 ;
        RECT 57.405 72.305 57.865 72.535 ;
        RECT 58.195 72.305 58.655 72.535 ;
        RECT 58.985 72.305 59.445 72.535 ;
        RECT 59.775 72.305 60.235 72.535 ;
        RECT 60.565 72.305 61.025 72.535 ;
        RECT 61.355 72.305 61.815 72.535 ;
        RECT 62.145 72.305 62.605 72.535 ;
        RECT 64.835 72.305 65.295 72.535 ;
        RECT 65.625 72.305 66.085 72.535 ;
        RECT 66.415 72.305 66.875 72.535 ;
        RECT 67.205 72.305 67.665 72.535 ;
        RECT 67.995 72.305 68.455 72.535 ;
        RECT 68.785 72.305 69.245 72.535 ;
        RECT 69.575 72.305 70.035 72.535 ;
        RECT 70.365 72.305 70.825 72.535 ;
        RECT 71.155 72.305 71.615 72.535 ;
        RECT 71.945 72.305 72.405 72.535 ;
        RECT 18.405 69.980 18.835 70.470 ;
        RECT 21.475 69.980 21.905 70.470 ;
        RECT 18.495 69.870 18.725 69.980 ;
        RECT 21.575 69.870 21.805 69.980 ;
        RECT 17.985 68.865 19.245 69.660 ;
        RECT 16.085 67.980 19.245 68.865 ;
        RECT 19.905 69.050 20.395 69.080 ;
        RECT 21.065 69.050 22.325 69.660 ;
        RECT 25.495 69.295 25.955 69.525 ;
        RECT 26.285 69.295 26.745 69.525 ;
        RECT 27.075 69.295 27.535 69.525 ;
        RECT 27.865 69.295 28.325 69.525 ;
        RECT 28.655 69.295 29.115 69.525 ;
        RECT 29.445 69.295 29.905 69.525 ;
        RECT 30.235 69.295 30.695 69.525 ;
        RECT 31.025 69.295 31.485 69.525 ;
        RECT 31.815 69.295 32.275 69.525 ;
        RECT 32.605 69.295 33.065 69.525 ;
        RECT 35.435 69.295 35.895 69.525 ;
        RECT 36.225 69.295 36.685 69.525 ;
        RECT 37.015 69.295 37.475 69.525 ;
        RECT 37.805 69.295 38.265 69.525 ;
        RECT 38.595 69.295 39.055 69.525 ;
        RECT 39.385 69.295 39.845 69.525 ;
        RECT 40.175 69.295 40.635 69.525 ;
        RECT 40.965 69.295 41.425 69.525 ;
        RECT 41.755 69.295 42.215 69.525 ;
        RECT 42.545 69.295 43.005 69.525 ;
        RECT 45.235 69.295 45.695 69.525 ;
        RECT 46.025 69.295 46.485 69.525 ;
        RECT 46.815 69.295 47.275 69.525 ;
        RECT 47.605 69.295 48.065 69.525 ;
        RECT 48.395 69.295 48.855 69.525 ;
        RECT 49.185 69.295 49.645 69.525 ;
        RECT 49.975 69.295 50.435 69.525 ;
        RECT 50.765 69.295 51.225 69.525 ;
        RECT 51.555 69.295 52.015 69.525 ;
        RECT 52.345 69.295 52.805 69.525 ;
        RECT 55.035 69.295 55.495 69.525 ;
        RECT 55.825 69.295 56.285 69.525 ;
        RECT 56.615 69.295 57.075 69.525 ;
        RECT 57.405 69.295 57.865 69.525 ;
        RECT 58.195 69.295 58.655 69.525 ;
        RECT 58.985 69.295 59.445 69.525 ;
        RECT 59.775 69.295 60.235 69.525 ;
        RECT 60.565 69.295 61.025 69.525 ;
        RECT 61.355 69.295 61.815 69.525 ;
        RECT 62.145 69.295 62.605 69.525 ;
        RECT 64.835 69.295 65.295 69.525 ;
        RECT 65.625 69.295 66.085 69.525 ;
        RECT 66.415 69.295 66.875 69.525 ;
        RECT 67.205 69.295 67.665 69.525 ;
        RECT 67.995 69.295 68.455 69.525 ;
        RECT 68.785 69.295 69.245 69.525 ;
        RECT 69.575 69.295 70.035 69.525 ;
        RECT 70.365 69.295 70.825 69.525 ;
        RECT 71.155 69.295 71.615 69.525 ;
        RECT 71.945 69.295 72.405 69.525 ;
        RECT 19.905 68.820 22.325 69.050 ;
        RECT 19.905 68.720 24.040 68.820 ;
        RECT 19.905 68.690 20.395 68.720 ;
        RECT 21.065 68.020 24.040 68.720 ;
        RECT 19.905 67.980 20.395 68.010 ;
        RECT 16.085 67.915 20.395 67.980 ;
        RECT 17.985 67.650 20.395 67.915 ;
        RECT 17.985 67.000 19.245 67.650 ;
        RECT 19.905 67.620 20.395 67.650 ;
        RECT 21.065 67.000 22.325 68.020 ;
        RECT 18.405 66.370 18.835 66.860 ;
        RECT 21.475 66.370 21.905 66.860 ;
        RECT 2.985 62.365 3.345 62.755 ;
        RECT 3.945 62.365 4.305 62.755 ;
        RECT 4.915 62.365 5.275 62.755 ;
        RECT 5.875 62.365 6.235 62.755 ;
        RECT 6.835 62.365 7.195 62.755 ;
        RECT 8.935 62.365 9.295 62.755 ;
        RECT 9.895 62.365 10.255 62.755 ;
        RECT 10.855 62.365 11.215 62.755 ;
        RECT 11.815 62.365 12.175 62.755 ;
        RECT 12.775 62.365 13.135 62.755 ;
        RECT 3.075 60.750 3.305 62.365 ;
        RECT 4.035 60.750 4.265 62.365 ;
        RECT 4.995 60.750 5.225 62.365 ;
        RECT 5.945 60.750 6.175 62.365 ;
        RECT 6.905 60.750 7.135 62.365 ;
        RECT 9.005 60.750 9.235 62.365 ;
        RECT 9.965 60.750 10.195 62.365 ;
        RECT 10.925 60.750 11.155 62.365 ;
        RECT 11.875 60.750 12.105 62.365 ;
        RECT 12.835 60.750 13.065 62.365 ;
        RECT 18.495 61.840 18.725 66.370 ;
        RECT 21.575 61.840 21.805 66.370 ;
        RECT 17.985 61.450 18.445 61.680 ;
        RECT 18.775 61.450 19.235 61.680 ;
        RECT 21.065 61.450 21.525 61.680 ;
        RECT 21.855 61.450 22.315 61.680 ;
        RECT 23.240 60.660 24.040 68.020 ;
        RECT 19.750 59.860 24.040 60.660 ;
        RECT 19.750 59.780 20.550 59.860 ;
        RECT 13.980 58.980 20.550 59.780 ;
        RECT 13.980 47.910 14.780 58.980 ;
        RECT 23.875 58.975 72.400 58.990 ;
        RECT 23.875 58.745 72.405 58.975 ;
        RECT 15.305 58.230 15.765 58.460 ;
        RECT 16.095 58.230 16.555 58.460 ;
        RECT 16.885 58.230 17.345 58.460 ;
        RECT 17.675 58.230 18.135 58.460 ;
        RECT 18.465 58.230 18.925 58.460 ;
        RECT 19.255 58.230 19.715 58.460 ;
        RECT 20.045 58.230 20.505 58.460 ;
        RECT 20.835 58.230 21.295 58.460 ;
        RECT 21.625 58.230 22.085 58.460 ;
        RECT 22.415 58.230 22.875 58.460 ;
        RECT 23.875 58.445 72.400 58.745 ;
        RECT 23.875 58.220 72.405 58.445 ;
        RECT 15.815 49.240 16.045 58.070 ;
        RECT 17.395 49.240 17.625 58.070 ;
        RECT 18.975 49.250 19.205 58.070 ;
        RECT 20.555 49.250 20.785 58.070 ;
        RECT 22.135 49.260 22.365 58.070 ;
        RECT 15.730 48.590 16.130 49.240 ;
        RECT 17.300 48.590 17.700 49.240 ;
        RECT 18.880 48.600 19.280 49.250 ;
        RECT 20.470 48.600 20.870 49.250 ;
        RECT 22.060 48.610 22.460 49.260 ;
        RECT 15.815 48.070 16.045 48.590 ;
        RECT 17.395 48.070 17.625 48.590 ;
        RECT 18.975 48.070 19.205 48.600 ;
        RECT 20.555 48.070 20.785 48.600 ;
        RECT 22.135 48.070 22.365 48.610 ;
        RECT 13.980 47.630 22.880 47.910 ;
        RECT 13.980 46.960 22.870 47.630 ;
        RECT 13.980 39.220 14.780 46.960 ;
        RECT 16.860 45.720 17.320 45.950 ;
        RECT 19.555 45.720 20.015 45.950 ;
        RECT 20.345 45.720 20.805 45.950 ;
        RECT 21.135 45.720 21.595 45.950 ;
        RECT 21.925 45.720 22.385 45.950 ;
        RECT 17.370 43.335 17.600 45.560 ;
        RECT 17.370 42.885 18.645 43.335 ;
        RECT 17.370 41.560 17.600 42.885 ;
        RECT 13.960 38.200 14.780 39.220 ;
        RECT 13.980 12.470 14.780 38.200 ;
        RECT 15.430 41.400 17.310 41.410 ;
        RECT 15.430 41.170 17.320 41.400 ;
        RECT 15.430 41.150 17.310 41.170 ;
        RECT 15.430 38.700 15.690 41.150 ;
        RECT 18.195 39.745 18.645 42.885 ;
        RECT 20.065 41.740 20.295 45.560 ;
        RECT 21.645 41.740 21.875 45.560 ;
        RECT 19.970 41.090 20.370 41.740 ;
        RECT 21.560 41.090 21.960 41.740 ;
        RECT 20.065 40.560 20.295 41.090 ;
        RECT 21.645 40.560 21.875 41.090 ;
        RECT 19.520 40.140 22.390 40.420 ;
        RECT 20.410 39.745 20.860 40.140 ;
        RECT 16.860 39.230 17.320 39.460 ;
        RECT 18.195 39.295 20.860 39.745 ;
        RECT 16.580 38.700 16.810 39.070 ;
        RECT 15.430 38.440 16.810 38.700 ;
        RECT 15.430 31.560 15.690 38.440 ;
        RECT 16.580 38.070 16.810 38.440 ;
        RECT 16.850 35.210 17.390 37.920 ;
        RECT 20.410 36.930 20.860 39.295 ;
        RECT 20.210 36.320 20.860 36.930 ;
        RECT 20.410 35.710 20.860 36.320 ;
        RECT 20.030 35.430 22.900 35.710 ;
        RECT 16.820 34.670 17.420 35.210 ;
        RECT 20.555 34.860 20.785 35.245 ;
        RECT 16.850 33.250 17.390 34.670 ;
        RECT 20.470 34.210 20.870 34.860 ;
        RECT 22.135 34.850 22.365 35.245 ;
        RECT 16.555 33.020 17.805 33.250 ;
        RECT 16.275 32.620 16.505 32.810 ;
        RECT 17.855 32.630 18.085 32.810 ;
        RECT 16.170 31.970 16.570 32.620 ;
        RECT 17.760 31.980 18.160 32.630 ;
        RECT 16.240 31.810 16.505 31.970 ;
        RECT 17.820 31.810 18.085 31.980 ;
        RECT 16.240 31.560 16.500 31.810 ;
        RECT 17.820 31.560 18.080 31.810 ;
        RECT 15.430 31.300 18.080 31.560 ;
        RECT 15.430 29.710 15.690 31.300 ;
        RECT 15.430 29.450 17.880 29.710 ;
        RECT 17.070 28.900 17.300 29.250 ;
        RECT 16.980 28.250 17.380 28.900 ;
        RECT 17.070 25.250 17.300 28.250 ;
        RECT 20.555 25.245 20.785 34.210 ;
        RECT 22.070 34.200 22.470 34.850 ;
        RECT 23.875 34.830 24.645 58.220 ;
        RECT 25.495 58.215 25.955 58.220 ;
        RECT 26.285 58.215 26.745 58.220 ;
        RECT 27.075 58.215 27.535 58.220 ;
        RECT 27.865 58.215 28.325 58.220 ;
        RECT 28.655 58.215 29.115 58.220 ;
        RECT 29.445 58.215 29.905 58.220 ;
        RECT 30.235 58.215 30.695 58.220 ;
        RECT 31.025 58.215 31.485 58.220 ;
        RECT 31.815 58.215 32.275 58.220 ;
        RECT 32.605 58.215 33.065 58.220 ;
        RECT 35.435 58.215 35.895 58.220 ;
        RECT 36.225 58.215 36.685 58.220 ;
        RECT 37.015 58.215 37.475 58.220 ;
        RECT 37.805 58.215 38.265 58.220 ;
        RECT 38.595 58.215 39.055 58.220 ;
        RECT 39.385 58.215 39.845 58.220 ;
        RECT 40.175 58.215 40.635 58.220 ;
        RECT 40.965 58.215 41.425 58.220 ;
        RECT 41.755 58.215 42.215 58.220 ;
        RECT 42.545 58.215 43.005 58.220 ;
        RECT 45.235 58.215 45.695 58.220 ;
        RECT 46.025 58.215 46.485 58.220 ;
        RECT 46.815 58.215 47.275 58.220 ;
        RECT 47.605 58.215 48.065 58.220 ;
        RECT 48.395 58.215 48.855 58.220 ;
        RECT 49.185 58.215 49.645 58.220 ;
        RECT 49.975 58.215 50.435 58.220 ;
        RECT 50.765 58.215 51.225 58.220 ;
        RECT 51.555 58.215 52.015 58.220 ;
        RECT 52.345 58.215 52.805 58.220 ;
        RECT 55.035 58.215 55.495 58.220 ;
        RECT 55.825 58.215 56.285 58.220 ;
        RECT 56.615 58.215 57.075 58.220 ;
        RECT 57.405 58.215 57.865 58.220 ;
        RECT 58.195 58.215 58.655 58.220 ;
        RECT 58.985 58.215 59.445 58.220 ;
        RECT 59.775 58.215 60.235 58.220 ;
        RECT 60.565 58.215 61.025 58.220 ;
        RECT 61.355 58.215 61.815 58.220 ;
        RECT 62.145 58.215 62.605 58.220 ;
        RECT 64.835 58.215 65.295 58.220 ;
        RECT 65.625 58.215 66.085 58.220 ;
        RECT 66.415 58.215 66.875 58.220 ;
        RECT 67.205 58.215 67.665 58.220 ;
        RECT 67.995 58.215 68.455 58.220 ;
        RECT 68.785 58.215 69.245 58.220 ;
        RECT 69.575 58.215 70.035 58.220 ;
        RECT 70.365 58.215 70.825 58.220 ;
        RECT 71.155 58.215 71.615 58.220 ;
        RECT 71.945 58.215 72.405 58.220 ;
        RECT 25.495 47.665 25.955 47.895 ;
        RECT 26.285 47.665 26.745 47.895 ;
        RECT 27.075 47.665 27.535 47.895 ;
        RECT 27.865 47.665 28.325 47.895 ;
        RECT 28.655 47.665 29.115 47.895 ;
        RECT 29.445 47.665 29.905 47.895 ;
        RECT 30.235 47.665 30.695 47.895 ;
        RECT 31.025 47.665 31.485 47.895 ;
        RECT 31.815 47.665 32.275 47.895 ;
        RECT 32.605 47.665 33.065 47.895 ;
        RECT 35.435 47.665 35.895 47.895 ;
        RECT 36.225 47.665 36.685 47.895 ;
        RECT 37.015 47.665 37.475 47.895 ;
        RECT 37.805 47.665 38.265 47.895 ;
        RECT 38.595 47.665 39.055 47.895 ;
        RECT 39.385 47.665 39.845 47.895 ;
        RECT 40.175 47.665 40.635 47.895 ;
        RECT 40.965 47.665 41.425 47.895 ;
        RECT 41.755 47.665 42.215 47.895 ;
        RECT 42.545 47.665 43.005 47.895 ;
        RECT 45.235 47.665 45.695 47.895 ;
        RECT 46.025 47.665 46.485 47.895 ;
        RECT 46.815 47.665 47.275 47.895 ;
        RECT 47.605 47.665 48.065 47.895 ;
        RECT 48.395 47.665 48.855 47.895 ;
        RECT 49.185 47.665 49.645 47.895 ;
        RECT 49.975 47.665 50.435 47.895 ;
        RECT 50.765 47.665 51.225 47.895 ;
        RECT 51.555 47.665 52.015 47.895 ;
        RECT 52.345 47.665 52.805 47.895 ;
        RECT 55.035 47.665 55.495 47.895 ;
        RECT 55.825 47.665 56.285 47.895 ;
        RECT 56.615 47.665 57.075 47.895 ;
        RECT 57.405 47.665 57.865 47.895 ;
        RECT 58.195 47.665 58.655 47.895 ;
        RECT 58.985 47.665 59.445 47.895 ;
        RECT 59.775 47.665 60.235 47.895 ;
        RECT 60.565 47.665 61.025 47.895 ;
        RECT 61.355 47.665 61.815 47.895 ;
        RECT 62.145 47.665 62.605 47.895 ;
        RECT 64.835 47.665 65.295 47.895 ;
        RECT 65.625 47.665 66.085 47.895 ;
        RECT 66.415 47.665 66.875 47.895 ;
        RECT 67.205 47.665 67.665 47.895 ;
        RECT 67.995 47.665 68.455 47.895 ;
        RECT 68.785 47.665 69.245 47.895 ;
        RECT 69.575 47.665 70.035 47.895 ;
        RECT 70.365 47.665 70.825 47.895 ;
        RECT 71.155 47.665 71.615 47.895 ;
        RECT 71.945 47.665 72.405 47.895 ;
        RECT 25.490 45.230 25.950 45.460 ;
        RECT 26.280 45.230 26.740 45.460 ;
        RECT 27.070 45.230 27.530 45.460 ;
        RECT 27.860 45.230 28.320 45.460 ;
        RECT 28.650 45.230 29.110 45.460 ;
        RECT 29.440 45.230 29.900 45.460 ;
        RECT 30.230 45.230 30.690 45.460 ;
        RECT 31.020 45.230 31.480 45.460 ;
        RECT 31.810 45.230 32.270 45.460 ;
        RECT 32.600 45.230 33.060 45.460 ;
        RECT 35.430 45.230 35.890 45.460 ;
        RECT 36.220 45.230 36.680 45.460 ;
        RECT 37.010 45.230 37.470 45.460 ;
        RECT 37.800 45.230 38.260 45.460 ;
        RECT 38.590 45.230 39.050 45.460 ;
        RECT 39.380 45.230 39.840 45.460 ;
        RECT 40.170 45.230 40.630 45.460 ;
        RECT 40.960 45.230 41.420 45.460 ;
        RECT 41.750 45.230 42.210 45.460 ;
        RECT 42.540 45.230 43.000 45.460 ;
        RECT 45.230 45.230 45.690 45.460 ;
        RECT 46.020 45.230 46.480 45.460 ;
        RECT 46.810 45.230 47.270 45.460 ;
        RECT 47.600 45.230 48.060 45.460 ;
        RECT 48.390 45.230 48.850 45.460 ;
        RECT 49.180 45.230 49.640 45.460 ;
        RECT 49.970 45.230 50.430 45.460 ;
        RECT 50.760 45.230 51.220 45.460 ;
        RECT 51.550 45.230 52.010 45.460 ;
        RECT 52.340 45.230 52.800 45.460 ;
        RECT 55.030 45.230 55.490 45.460 ;
        RECT 55.820 45.230 56.280 45.460 ;
        RECT 56.610 45.230 57.070 45.460 ;
        RECT 57.400 45.230 57.860 45.460 ;
        RECT 58.190 45.230 58.650 45.460 ;
        RECT 58.980 45.230 59.440 45.460 ;
        RECT 59.770 45.230 60.230 45.460 ;
        RECT 60.560 45.230 61.020 45.460 ;
        RECT 61.350 45.230 61.810 45.460 ;
        RECT 62.140 45.230 62.600 45.460 ;
        RECT 64.830 45.230 65.290 45.460 ;
        RECT 65.620 45.230 66.080 45.460 ;
        RECT 66.410 45.230 66.870 45.460 ;
        RECT 67.200 45.230 67.660 45.460 ;
        RECT 67.990 45.230 68.450 45.460 ;
        RECT 68.780 45.230 69.240 45.460 ;
        RECT 69.570 45.230 70.030 45.460 ;
        RECT 70.360 45.230 70.820 45.460 ;
        RECT 71.150 45.230 71.610 45.460 ;
        RECT 71.940 45.230 72.400 45.460 ;
        RECT 22.135 25.245 22.365 34.200 ;
        RECT 23.875 34.060 72.400 34.830 ;
        RECT 16.560 24.810 17.020 25.040 ;
        RECT 17.350 24.810 17.810 25.040 ;
        RECT 20.045 24.805 20.505 25.035 ;
        RECT 20.835 24.805 21.295 25.035 ;
        RECT 21.625 24.805 22.085 25.035 ;
        RECT 22.415 24.805 22.875 25.035 ;
        RECT 15.305 22.875 15.765 23.105 ;
        RECT 16.095 22.875 16.555 23.105 ;
        RECT 16.885 22.875 17.345 23.105 ;
        RECT 17.675 22.875 18.135 23.105 ;
        RECT 18.465 22.875 18.925 23.105 ;
        RECT 19.255 22.875 19.715 23.105 ;
        RECT 20.045 22.875 20.505 23.105 ;
        RECT 20.835 22.875 21.295 23.105 ;
        RECT 21.625 22.875 22.085 23.105 ;
        RECT 22.415 22.875 22.875 23.105 ;
        RECT 15.815 13.810 16.045 22.665 ;
        RECT 15.730 13.160 16.130 13.810 ;
        RECT 17.395 13.800 17.625 22.665 ;
        RECT 18.975 13.800 19.205 22.665 ;
        RECT 15.815 12.665 16.045 13.160 ;
        RECT 17.310 13.150 17.710 13.800 ;
        RECT 18.880 13.150 19.280 13.800 ;
        RECT 20.555 13.790 20.785 22.665 ;
        RECT 22.135 13.790 22.365 22.665 ;
        RECT 17.395 12.665 17.625 13.150 ;
        RECT 18.975 12.665 19.205 13.150 ;
        RECT 20.460 13.140 20.860 13.790 ;
        RECT 22.030 13.140 22.430 13.790 ;
        RECT 23.875 13.360 24.645 34.060 ;
        RECT 25.490 34.050 25.950 34.060 ;
        RECT 26.280 34.050 26.740 34.060 ;
        RECT 27.070 34.050 27.530 34.060 ;
        RECT 27.860 34.050 28.320 34.060 ;
        RECT 28.650 34.050 29.110 34.060 ;
        RECT 29.440 34.050 29.900 34.060 ;
        RECT 30.230 34.050 30.690 34.060 ;
        RECT 31.020 34.050 31.480 34.060 ;
        RECT 31.810 34.050 32.270 34.060 ;
        RECT 32.600 34.050 33.060 34.060 ;
        RECT 35.430 34.050 35.890 34.060 ;
        RECT 36.220 34.050 36.680 34.060 ;
        RECT 37.010 34.050 37.470 34.060 ;
        RECT 37.800 34.050 38.260 34.060 ;
        RECT 38.590 34.050 39.050 34.060 ;
        RECT 39.380 34.050 39.840 34.060 ;
        RECT 40.170 34.050 40.630 34.060 ;
        RECT 40.960 34.050 41.420 34.060 ;
        RECT 41.750 34.050 42.210 34.060 ;
        RECT 42.540 34.050 43.000 34.060 ;
        RECT 45.230 34.050 45.690 34.060 ;
        RECT 46.020 34.050 46.480 34.060 ;
        RECT 46.810 34.050 47.270 34.060 ;
        RECT 47.600 34.050 48.060 34.060 ;
        RECT 48.390 34.050 48.850 34.060 ;
        RECT 49.180 34.050 49.640 34.060 ;
        RECT 49.970 34.050 50.430 34.060 ;
        RECT 50.760 34.050 51.220 34.060 ;
        RECT 51.550 34.050 52.010 34.060 ;
        RECT 52.340 34.050 52.800 34.060 ;
        RECT 55.030 34.050 55.490 34.060 ;
        RECT 55.820 34.050 56.280 34.060 ;
        RECT 56.610 34.050 57.070 34.060 ;
        RECT 57.400 34.050 57.860 34.060 ;
        RECT 58.190 34.050 58.650 34.060 ;
        RECT 58.980 34.050 59.440 34.060 ;
        RECT 59.770 34.050 60.230 34.060 ;
        RECT 60.560 34.050 61.020 34.060 ;
        RECT 61.350 34.050 61.810 34.060 ;
        RECT 62.140 34.050 62.600 34.060 ;
        RECT 64.830 34.050 65.290 34.060 ;
        RECT 65.620 34.050 66.080 34.060 ;
        RECT 66.410 34.050 66.870 34.060 ;
        RECT 67.200 34.050 67.660 34.060 ;
        RECT 67.990 34.050 68.450 34.060 ;
        RECT 68.780 34.050 69.240 34.060 ;
        RECT 69.570 34.050 70.030 34.060 ;
        RECT 70.360 34.050 70.820 34.060 ;
        RECT 71.150 34.050 71.610 34.060 ;
        RECT 71.940 34.050 72.400 34.060 ;
        RECT 25.490 23.410 25.950 23.640 ;
        RECT 26.280 23.410 26.740 23.640 ;
        RECT 27.070 23.410 27.530 23.640 ;
        RECT 27.860 23.410 28.320 23.640 ;
        RECT 28.650 23.410 29.110 23.640 ;
        RECT 29.440 23.410 29.900 23.640 ;
        RECT 30.230 23.410 30.690 23.640 ;
        RECT 31.020 23.410 31.480 23.640 ;
        RECT 31.810 23.410 32.270 23.640 ;
        RECT 32.600 23.410 33.060 23.640 ;
        RECT 35.430 23.410 35.890 23.640 ;
        RECT 36.220 23.410 36.680 23.640 ;
        RECT 37.010 23.410 37.470 23.640 ;
        RECT 37.800 23.410 38.260 23.640 ;
        RECT 38.590 23.410 39.050 23.640 ;
        RECT 39.380 23.410 39.840 23.640 ;
        RECT 40.170 23.410 40.630 23.640 ;
        RECT 40.960 23.410 41.420 23.640 ;
        RECT 41.750 23.410 42.210 23.640 ;
        RECT 42.540 23.410 43.000 23.640 ;
        RECT 45.230 23.410 45.690 23.640 ;
        RECT 46.020 23.410 46.480 23.640 ;
        RECT 46.810 23.410 47.270 23.640 ;
        RECT 47.600 23.410 48.060 23.640 ;
        RECT 48.390 23.410 48.850 23.640 ;
        RECT 49.180 23.410 49.640 23.640 ;
        RECT 49.970 23.410 50.430 23.640 ;
        RECT 50.760 23.410 51.220 23.640 ;
        RECT 51.550 23.410 52.010 23.640 ;
        RECT 52.340 23.410 52.800 23.640 ;
        RECT 55.030 23.410 55.490 23.640 ;
        RECT 55.820 23.410 56.280 23.640 ;
        RECT 56.610 23.410 57.070 23.640 ;
        RECT 57.400 23.410 57.860 23.640 ;
        RECT 58.190 23.410 58.650 23.640 ;
        RECT 58.980 23.410 59.440 23.640 ;
        RECT 59.770 23.410 60.230 23.640 ;
        RECT 60.560 23.410 61.020 23.640 ;
        RECT 61.350 23.410 61.810 23.640 ;
        RECT 62.140 23.410 62.600 23.640 ;
        RECT 64.830 23.410 65.290 23.640 ;
        RECT 65.620 23.410 66.080 23.640 ;
        RECT 66.410 23.410 66.870 23.640 ;
        RECT 67.200 23.410 67.660 23.640 ;
        RECT 67.990 23.410 68.450 23.640 ;
        RECT 68.780 23.410 69.240 23.640 ;
        RECT 69.570 23.410 70.030 23.640 ;
        RECT 70.360 23.410 70.820 23.640 ;
        RECT 71.150 23.410 71.610 23.640 ;
        RECT 71.940 23.410 72.400 23.640 ;
        RECT 25.490 22.870 25.950 23.100 ;
        RECT 26.280 22.870 26.740 23.100 ;
        RECT 27.070 22.870 27.530 23.100 ;
        RECT 27.860 22.870 28.320 23.100 ;
        RECT 28.650 22.870 29.110 23.100 ;
        RECT 29.440 22.870 29.900 23.100 ;
        RECT 30.230 22.870 30.690 23.100 ;
        RECT 31.020 22.870 31.480 23.100 ;
        RECT 31.810 22.870 32.270 23.100 ;
        RECT 32.600 22.870 33.060 23.100 ;
        RECT 35.430 22.870 35.890 23.100 ;
        RECT 36.220 22.870 36.680 23.100 ;
        RECT 37.010 22.870 37.470 23.100 ;
        RECT 37.800 22.870 38.260 23.100 ;
        RECT 38.590 22.870 39.050 23.100 ;
        RECT 39.380 22.870 39.840 23.100 ;
        RECT 40.170 22.870 40.630 23.100 ;
        RECT 40.960 22.870 41.420 23.100 ;
        RECT 41.750 22.870 42.210 23.100 ;
        RECT 42.540 22.870 43.000 23.100 ;
        RECT 45.230 22.870 45.690 23.100 ;
        RECT 46.020 22.870 46.480 23.100 ;
        RECT 46.810 22.870 47.270 23.100 ;
        RECT 47.600 22.870 48.060 23.100 ;
        RECT 48.390 22.870 48.850 23.100 ;
        RECT 49.180 22.870 49.640 23.100 ;
        RECT 49.970 22.870 50.430 23.100 ;
        RECT 50.760 22.870 51.220 23.100 ;
        RECT 51.550 22.870 52.010 23.100 ;
        RECT 52.340 22.870 52.800 23.100 ;
        RECT 55.030 22.870 55.490 23.100 ;
        RECT 55.820 22.870 56.280 23.100 ;
        RECT 56.610 22.870 57.070 23.100 ;
        RECT 57.400 22.870 57.860 23.100 ;
        RECT 58.190 22.870 58.650 23.100 ;
        RECT 58.980 22.870 59.440 23.100 ;
        RECT 59.770 22.870 60.230 23.100 ;
        RECT 60.560 22.870 61.020 23.100 ;
        RECT 61.350 22.870 61.810 23.100 ;
        RECT 62.140 22.870 62.600 23.100 ;
        RECT 64.830 22.870 65.290 23.100 ;
        RECT 65.620 22.870 66.080 23.100 ;
        RECT 66.410 22.870 66.870 23.100 ;
        RECT 67.200 22.870 67.660 23.100 ;
        RECT 67.990 22.870 68.450 23.100 ;
        RECT 68.780 22.870 69.240 23.100 ;
        RECT 69.570 22.870 70.030 23.100 ;
        RECT 70.360 22.870 70.820 23.100 ;
        RECT 71.150 22.870 71.610 23.100 ;
        RECT 71.940 22.870 72.400 23.100 ;
        RECT 20.555 12.665 20.785 13.140 ;
        RECT 22.135 12.665 22.365 13.140 ;
        RECT 23.860 12.475 24.660 13.360 ;
        RECT 23.860 12.470 26.215 12.475 ;
        RECT 13.980 11.670 22.900 12.470 ;
        RECT 23.860 11.750 72.400 12.470 ;
        RECT 23.875 11.705 72.400 11.750 ;
        RECT 25.490 11.690 25.950 11.705 ;
        RECT 26.215 11.700 72.400 11.705 ;
        RECT 26.280 11.690 26.740 11.700 ;
        RECT 27.070 11.690 27.530 11.700 ;
        RECT 27.860 11.690 28.320 11.700 ;
        RECT 28.650 11.690 29.110 11.700 ;
        RECT 29.440 11.690 29.900 11.700 ;
        RECT 30.230 11.690 30.690 11.700 ;
        RECT 31.020 11.690 31.480 11.700 ;
        RECT 31.810 11.690 32.270 11.700 ;
        RECT 32.600 11.690 33.060 11.700 ;
        RECT 35.430 11.690 35.890 11.700 ;
        RECT 36.220 11.690 36.680 11.700 ;
        RECT 37.010 11.690 37.470 11.700 ;
        RECT 37.800 11.690 38.260 11.700 ;
        RECT 38.590 11.690 39.050 11.700 ;
        RECT 39.380 11.690 39.840 11.700 ;
        RECT 40.170 11.690 40.630 11.700 ;
        RECT 40.960 11.690 41.420 11.700 ;
        RECT 41.750 11.690 42.210 11.700 ;
        RECT 42.540 11.690 43.000 11.700 ;
        RECT 45.230 11.690 45.690 11.700 ;
        RECT 46.020 11.690 46.480 11.700 ;
        RECT 46.810 11.690 47.270 11.700 ;
        RECT 47.600 11.690 48.060 11.700 ;
        RECT 48.390 11.690 48.850 11.700 ;
        RECT 49.180 11.690 49.640 11.700 ;
        RECT 49.970 11.690 50.430 11.700 ;
        RECT 50.760 11.690 51.220 11.700 ;
        RECT 51.550 11.690 52.010 11.700 ;
        RECT 52.340 11.690 52.800 11.700 ;
        RECT 55.030 11.690 55.490 11.700 ;
        RECT 55.820 11.690 56.280 11.700 ;
        RECT 56.610 11.690 57.070 11.700 ;
        RECT 57.400 11.690 57.860 11.700 ;
        RECT 58.190 11.690 58.650 11.700 ;
        RECT 58.980 11.690 59.440 11.700 ;
        RECT 59.770 11.690 60.230 11.700 ;
        RECT 60.560 11.690 61.020 11.700 ;
        RECT 61.350 11.690 61.810 11.700 ;
        RECT 62.140 11.690 62.600 11.700 ;
        RECT 64.830 11.690 65.290 11.700 ;
        RECT 65.620 11.690 66.080 11.700 ;
        RECT 66.410 11.690 66.870 11.700 ;
        RECT 67.200 11.690 67.660 11.700 ;
        RECT 67.990 11.690 68.450 11.700 ;
        RECT 68.780 11.690 69.240 11.700 ;
        RECT 69.570 11.690 70.030 11.700 ;
        RECT 70.360 11.690 70.820 11.700 ;
        RECT 71.150 11.690 71.610 11.700 ;
        RECT 71.940 11.690 72.400 11.700 ;
        RECT 15.815 11.120 16.045 11.485 ;
        RECT 17.395 11.120 17.625 11.485 ;
        RECT 18.975 11.120 19.215 11.485 ;
        RECT 20.555 11.130 20.785 11.485 ;
        RECT 22.135 11.130 22.365 11.485 ;
        RECT 15.720 10.470 16.120 11.120 ;
        RECT 17.310 10.470 17.710 11.120 ;
        RECT 18.890 10.470 19.290 11.120 ;
        RECT 20.450 10.480 20.850 11.130 ;
        RECT 22.030 10.480 22.430 11.130 ;
        RECT 15.815 1.485 16.045 10.470 ;
        RECT 17.395 1.485 17.625 10.470 ;
        RECT 18.975 1.485 19.215 10.470 ;
        RECT 20.555 1.485 20.785 10.480 ;
        RECT 22.135 1.485 22.365 10.480 ;
        RECT 15.305 1.045 15.765 1.275 ;
        RECT 16.095 1.045 16.555 1.275 ;
        RECT 16.885 1.045 17.345 1.275 ;
        RECT 17.675 1.045 18.135 1.275 ;
        RECT 18.465 1.045 18.925 1.275 ;
        RECT 19.255 1.045 19.715 1.275 ;
        RECT 20.045 1.045 20.505 1.275 ;
        RECT 20.835 1.045 21.295 1.275 ;
        RECT 21.625 1.045 22.085 1.275 ;
        RECT 22.415 1.045 22.875 1.275 ;
        RECT 25.490 1.050 25.950 1.280 ;
        RECT 26.280 1.050 26.740 1.280 ;
        RECT 27.070 1.050 27.530 1.280 ;
        RECT 27.860 1.050 28.320 1.280 ;
        RECT 28.650 1.050 29.110 1.280 ;
        RECT 29.440 1.050 29.900 1.280 ;
        RECT 30.230 1.050 30.690 1.280 ;
        RECT 31.020 1.050 31.480 1.280 ;
        RECT 31.810 1.050 32.270 1.280 ;
        RECT 32.600 1.050 33.060 1.280 ;
        RECT 35.430 1.050 35.890 1.280 ;
        RECT 36.220 1.050 36.680 1.280 ;
        RECT 37.010 1.050 37.470 1.280 ;
        RECT 37.800 1.050 38.260 1.280 ;
        RECT 38.590 1.050 39.050 1.280 ;
        RECT 39.380 1.050 39.840 1.280 ;
        RECT 40.170 1.050 40.630 1.280 ;
        RECT 40.960 1.050 41.420 1.280 ;
        RECT 41.750 1.050 42.210 1.280 ;
        RECT 42.540 1.050 43.000 1.280 ;
        RECT 45.230 1.050 45.690 1.280 ;
        RECT 46.020 1.050 46.480 1.280 ;
        RECT 46.810 1.050 47.270 1.280 ;
        RECT 47.600 1.050 48.060 1.280 ;
        RECT 48.390 1.050 48.850 1.280 ;
        RECT 49.180 1.050 49.640 1.280 ;
        RECT 49.970 1.050 50.430 1.280 ;
        RECT 50.760 1.050 51.220 1.280 ;
        RECT 51.550 1.050 52.010 1.280 ;
        RECT 52.340 1.050 52.800 1.280 ;
        RECT 55.030 1.050 55.490 1.280 ;
        RECT 55.820 1.050 56.280 1.280 ;
        RECT 56.610 1.050 57.070 1.280 ;
        RECT 57.400 1.050 57.860 1.280 ;
        RECT 58.190 1.050 58.650 1.280 ;
        RECT 58.980 1.050 59.440 1.280 ;
        RECT 59.770 1.050 60.230 1.280 ;
        RECT 60.560 1.050 61.020 1.280 ;
        RECT 61.350 1.050 61.810 1.280 ;
        RECT 62.140 1.050 62.600 1.280 ;
        RECT 64.830 1.050 65.290 1.280 ;
        RECT 65.620 1.050 66.080 1.280 ;
        RECT 66.410 1.050 66.870 1.280 ;
        RECT 67.200 1.050 67.660 1.280 ;
        RECT 67.990 1.050 68.450 1.280 ;
        RECT 68.780 1.050 69.240 1.280 ;
        RECT 69.570 1.050 70.030 1.280 ;
        RECT 70.360 1.050 70.820 1.280 ;
        RECT 71.150 1.050 71.610 1.280 ;
        RECT 71.940 1.050 72.400 1.280 ;
      LAYER via ;
        RECT 15.770 130.710 16.070 131.360 ;
        RECT 17.360 130.710 17.660 131.360 ;
        RECT 18.940 130.710 19.240 131.360 ;
        RECT 20.500 130.700 20.800 131.350 ;
        RECT 22.080 130.700 22.380 131.350 ;
        RECT 15.780 128.020 16.080 128.670 ;
        RECT 17.360 128.030 17.660 128.680 ;
        RECT 18.930 128.030 19.230 128.680 ;
        RECT 20.510 128.040 20.810 128.690 ;
        RECT 22.080 128.040 22.380 128.690 ;
        RECT 23.910 128.470 24.610 130.080 ;
        RECT 17.030 112.930 17.330 113.580 ;
        RECT 14.010 102.610 14.710 103.630 ;
        RECT 16.220 109.210 16.520 109.860 ;
        RECT 17.810 109.200 18.110 109.850 ;
        RECT 20.520 106.970 20.820 107.620 ;
        RECT 22.120 106.980 22.420 107.630 ;
        RECT 16.850 106.390 17.390 106.930 ;
        RECT 20.260 104.900 20.800 105.510 ;
        RECT 20.020 100.090 20.320 100.740 ;
        RECT 21.610 100.090 21.910 100.740 ;
        RECT 4.095 78.455 4.385 79.055 ;
        RECT 5.675 78.455 5.965 79.055 ;
        RECT 7.255 78.455 7.545 79.055 ;
        RECT 8.595 78.455 8.885 79.055 ;
        RECT 10.175 78.455 10.465 79.055 ;
        RECT 11.755 78.455 12.045 79.055 ;
        RECT 15.780 92.590 16.080 93.240 ;
        RECT 17.350 92.590 17.650 93.240 ;
        RECT 18.930 92.580 19.230 93.230 ;
        RECT 20.520 92.580 20.820 93.230 ;
        RECT 22.110 92.570 22.410 93.220 ;
        RECT 23.950 92.360 24.560 93.650 ;
        RECT 8.935 77.605 9.195 77.865 ;
        RECT 0.945 73.615 1.255 74.775 ;
        RECT 3.335 73.615 3.645 74.775 ;
        RECT 2.165 65.315 2.425 65.705 ;
        RECT 5.715 73.615 6.025 74.775 ;
        RECT 4.545 65.315 4.805 65.705 ;
        RECT 9.995 73.615 10.305 74.775 ;
        RECT 6.925 65.315 7.185 65.705 ;
        RECT 8.825 65.315 9.085 65.705 ;
        RECT 12.375 73.615 12.685 74.775 ;
        RECT 11.205 65.315 11.465 65.705 ;
        RECT 14.755 73.615 15.065 74.775 ;
        RECT 13.585 65.315 13.845 65.705 ;
        RECT 18.455 69.980 18.785 70.470 ;
        RECT 21.525 69.980 21.855 70.470 ;
        RECT 19.905 67.650 20.395 67.980 ;
        RECT 18.455 66.370 18.785 66.860 ;
        RECT 21.525 66.370 21.855 66.860 ;
        RECT 3.035 62.365 3.295 62.755 ;
        RECT 3.995 62.365 4.255 62.755 ;
        RECT 4.965 62.365 5.225 62.755 ;
        RECT 5.925 62.365 6.185 62.755 ;
        RECT 6.885 62.365 7.145 62.755 ;
        RECT 8.985 62.365 9.245 62.755 ;
        RECT 9.945 62.365 10.205 62.755 ;
        RECT 10.905 62.365 11.165 62.755 ;
        RECT 11.865 62.365 12.125 62.755 ;
        RECT 12.825 62.365 13.085 62.755 ;
        RECT 15.780 48.590 16.080 49.240 ;
        RECT 17.350 48.590 17.650 49.240 ;
        RECT 18.930 48.600 19.230 49.250 ;
        RECT 20.520 48.600 20.820 49.250 ;
        RECT 22.110 48.610 22.410 49.260 ;
        RECT 23.950 48.180 24.560 49.470 ;
        RECT 14.010 38.200 14.710 39.220 ;
        RECT 20.020 41.090 20.320 41.740 ;
        RECT 21.610 41.090 21.910 41.740 ;
        RECT 20.260 36.320 20.800 36.930 ;
        RECT 16.850 34.670 17.390 35.210 ;
        RECT 20.520 34.210 20.820 34.860 ;
        RECT 16.220 31.970 16.520 32.620 ;
        RECT 17.810 31.980 18.110 32.630 ;
        RECT 17.030 28.250 17.330 28.900 ;
        RECT 22.120 34.200 22.420 34.850 ;
        RECT 15.780 13.160 16.080 13.810 ;
        RECT 17.360 13.150 17.660 13.800 ;
        RECT 18.930 13.150 19.230 13.800 ;
        RECT 20.510 13.140 20.810 13.790 ;
        RECT 22.080 13.140 22.380 13.790 ;
        RECT 23.910 11.750 24.610 13.360 ;
        RECT 15.770 10.470 16.070 11.120 ;
        RECT 17.360 10.470 17.660 11.120 ;
        RECT 18.940 10.470 19.240 11.120 ;
        RECT 20.500 10.480 20.800 11.130 ;
        RECT 22.080 10.480 22.380 11.130 ;
      LAYER met2 ;
        RECT 15.770 131.240 16.070 131.410 ;
        RECT 17.360 131.240 17.660 131.410 ;
        RECT 18.940 131.240 19.240 131.410 ;
        RECT 20.500 131.240 20.800 131.400 ;
        RECT 22.080 131.240 22.380 131.400 ;
        RECT 15.770 130.820 24.250 131.240 ;
        RECT 15.770 130.660 16.070 130.820 ;
        RECT 17.360 130.660 17.660 130.820 ;
        RECT 18.940 130.660 19.240 130.820 ;
        RECT 20.500 130.650 20.800 130.820 ;
        RECT 22.080 130.650 22.380 130.820 ;
        RECT 23.830 130.130 24.250 130.820 ;
        RECT 15.780 128.590 16.080 128.720 ;
        RECT 17.360 128.590 17.660 128.730 ;
        RECT 18.930 128.590 19.230 128.730 ;
        RECT 20.510 128.590 20.810 128.740 ;
        RECT 22.080 128.590 22.380 128.740 ;
        RECT 23.830 128.590 24.610 130.130 ;
        RECT 15.780 128.420 24.610 128.590 ;
        RECT 15.780 128.170 24.250 128.420 ;
        RECT 15.780 127.970 16.080 128.170 ;
        RECT 17.360 127.980 17.660 128.170 ;
        RECT 18.930 127.980 19.230 128.170 ;
        RECT 20.510 127.990 20.810 128.170 ;
        RECT 22.080 127.990 22.380 128.170 ;
        RECT 17.030 113.420 17.330 113.630 ;
        RECT 15.460 113.030 17.330 113.420 ;
        RECT 15.460 105.395 15.850 113.030 ;
        RECT 17.030 112.880 17.330 113.030 ;
        RECT 16.220 109.160 16.520 109.910 ;
        RECT 17.810 109.150 18.110 109.900 ;
        RECT 20.520 107.540 20.820 107.670 ;
        RECT 22.120 107.540 22.420 107.680 ;
        RECT 20.520 107.070 22.420 107.540 ;
        RECT 16.850 106.930 17.390 106.960 ;
        RECT 16.805 106.390 17.435 106.930 ;
        RECT 20.520 106.920 20.820 107.070 ;
        RECT 16.850 106.360 17.390 106.390 ;
        RECT 20.260 105.395 20.800 105.560 ;
        RECT 15.460 105.005 20.800 105.395 ;
        RECT 20.260 104.850 20.800 105.005 ;
        RECT 14.010 103.315 14.710 103.680 ;
        RECT 21.095 103.315 21.525 107.070 ;
        RECT 22.120 106.930 22.420 107.070 ;
        RECT 14.010 102.885 21.525 103.315 ;
        RECT 14.010 102.560 14.710 102.885 ;
        RECT 21.095 100.790 21.525 102.885 ;
        RECT 20.020 100.640 20.320 100.790 ;
        RECT 21.095 100.640 21.910 100.790 ;
        RECT 20.020 100.210 21.910 100.640 ;
        RECT 20.020 100.040 20.320 100.210 ;
        RECT 21.610 100.040 21.910 100.210 ;
        RECT 15.780 93.180 16.080 93.290 ;
        RECT 17.350 93.180 17.650 93.290 ;
        RECT 18.930 93.180 19.230 93.280 ;
        RECT 20.520 93.180 20.820 93.280 ;
        RECT 22.110 93.180 22.410 93.270 ;
        RECT 23.950 93.180 24.560 93.700 ;
        RECT 15.780 92.650 24.560 93.180 ;
        RECT 15.780 92.540 16.080 92.650 ;
        RECT 17.350 92.540 17.650 92.650 ;
        RECT 18.930 92.530 19.230 92.650 ;
        RECT 20.520 92.530 20.820 92.650 ;
        RECT 22.110 92.520 22.410 92.650 ;
        RECT 23.950 92.310 24.560 92.650 ;
        RECT 4.095 79.055 4.385 79.105 ;
        RECT 5.675 79.055 5.965 79.105 ;
        RECT 7.255 79.055 7.545 79.105 ;
        RECT 3.335 78.455 7.545 79.055 ;
        RECT 4.095 78.405 4.385 78.455 ;
        RECT 4.855 78.405 5.965 78.455 ;
        RECT 7.255 78.405 7.545 78.455 ;
        RECT 8.595 79.055 8.885 79.105 ;
        RECT 10.175 79.055 10.465 79.105 ;
        RECT 11.755 79.055 12.045 79.105 ;
        RECT 8.595 78.455 12.805 79.055 ;
        RECT 8.595 78.405 8.885 78.455 ;
        RECT 10.175 78.410 11.215 78.455 ;
        RECT 10.175 78.405 11.145 78.410 ;
        RECT 11.755 78.405 12.045 78.455 ;
        RECT 0.945 74.775 1.255 74.825 ;
        RECT 3.335 74.775 3.645 74.825 ;
        RECT 4.855 74.775 5.345 78.405 ;
        RECT 7.285 78.255 7.525 78.405 ;
        RECT 7.285 78.015 8.295 78.255 ;
        RECT 8.015 77.855 8.295 78.015 ;
        RECT 8.935 77.855 9.195 77.895 ;
        RECT 8.015 77.615 9.195 77.855 ;
        RECT 8.935 77.575 9.195 77.615 ;
        RECT 5.715 74.775 6.025 74.825 ;
        RECT 0.945 73.615 6.025 74.775 ;
        RECT 0.945 73.565 1.255 73.615 ;
        RECT 3.335 73.565 3.645 73.615 ;
        RECT 5.715 73.565 6.025 73.615 ;
        RECT 9.995 74.775 10.305 74.825 ;
        RECT 10.655 74.775 11.145 78.405 ;
        RECT 12.375 74.775 12.685 74.825 ;
        RECT 14.755 74.775 15.065 74.825 ;
        RECT 9.995 73.615 15.065 74.775 ;
        RECT 9.995 73.565 10.305 73.615 ;
        RECT 12.375 73.565 12.685 73.615 ;
        RECT 14.755 73.565 15.065 73.615 ;
        RECT 18.455 69.050 18.785 70.520 ;
        RECT 18.455 68.720 20.425 69.050 ;
        RECT 18.455 66.320 18.785 68.720 ;
        RECT 21.525 67.980 21.855 70.520 ;
        RECT 19.875 67.650 21.855 67.980 ;
        RECT 21.525 66.320 21.855 67.650 ;
        RECT 2.165 64.455 2.425 65.755 ;
        RECT 4.545 64.455 4.805 65.755 ;
        RECT 6.925 64.455 7.185 65.755 ;
        RECT 2.165 64.025 7.185 64.455 ;
        RECT 8.825 64.455 9.085 65.755 ;
        RECT 11.205 64.455 11.465 65.755 ;
        RECT 13.585 64.455 13.845 65.755 ;
        RECT 8.825 64.025 13.845 64.455 ;
        RECT 2.505 63.485 7.525 64.025 ;
        RECT 8.605 63.485 13.625 64.025 ;
        RECT 3.035 62.315 3.295 63.485 ;
        RECT 3.995 62.315 4.255 63.485 ;
        RECT 4.965 62.315 5.225 63.485 ;
        RECT 5.925 62.315 6.185 63.485 ;
        RECT 6.885 62.315 7.145 63.485 ;
        RECT 8.985 62.315 9.245 63.485 ;
        RECT 9.945 62.315 10.205 63.485 ;
        RECT 10.905 62.315 11.165 63.485 ;
        RECT 11.865 62.315 12.125 63.485 ;
        RECT 12.825 62.315 13.085 63.485 ;
        RECT 15.780 49.180 16.080 49.290 ;
        RECT 17.350 49.180 17.650 49.290 ;
        RECT 18.930 49.180 19.230 49.300 ;
        RECT 20.520 49.180 20.820 49.300 ;
        RECT 22.110 49.180 22.410 49.310 ;
        RECT 23.950 49.180 24.560 49.520 ;
        RECT 15.780 48.650 24.560 49.180 ;
        RECT 15.780 48.540 16.080 48.650 ;
        RECT 17.350 48.540 17.650 48.650 ;
        RECT 18.930 48.550 19.230 48.650 ;
        RECT 20.520 48.550 20.820 48.650 ;
        RECT 22.110 48.560 22.410 48.650 ;
        RECT 23.950 48.130 24.560 48.650 ;
        RECT 20.020 41.620 20.320 41.790 ;
        RECT 21.610 41.620 21.910 41.790 ;
        RECT 20.020 41.190 21.910 41.620 ;
        RECT 20.020 41.040 20.320 41.190 ;
        RECT 21.095 41.040 21.910 41.190 ;
        RECT 14.010 38.945 14.710 39.270 ;
        RECT 21.095 38.945 21.525 41.040 ;
        RECT 14.010 38.515 21.525 38.945 ;
        RECT 14.010 38.150 14.710 38.515 ;
        RECT 20.260 36.825 20.800 36.980 ;
        RECT 15.460 36.435 20.800 36.825 ;
        RECT 15.460 28.800 15.850 36.435 ;
        RECT 20.260 36.270 20.800 36.435 ;
        RECT 16.850 35.210 17.390 35.240 ;
        RECT 16.805 34.670 17.435 35.210 ;
        RECT 20.520 34.760 20.820 34.910 ;
        RECT 21.095 34.760 21.525 38.515 ;
        RECT 22.120 34.760 22.420 34.900 ;
        RECT 16.850 34.640 17.390 34.670 ;
        RECT 20.520 34.290 22.420 34.760 ;
        RECT 20.520 34.160 20.820 34.290 ;
        RECT 22.120 34.150 22.420 34.290 ;
        RECT 16.220 31.920 16.520 32.670 ;
        RECT 17.810 31.930 18.110 32.680 ;
        RECT 17.030 28.800 17.330 28.950 ;
        RECT 15.460 28.410 17.330 28.800 ;
        RECT 17.030 28.200 17.330 28.410 ;
        RECT 15.780 13.660 16.080 13.860 ;
        RECT 17.360 13.660 17.660 13.850 ;
        RECT 18.930 13.660 19.230 13.850 ;
        RECT 20.510 13.660 20.810 13.840 ;
        RECT 22.080 13.660 22.380 13.840 ;
        RECT 15.780 13.410 24.250 13.660 ;
        RECT 15.780 13.240 24.610 13.410 ;
        RECT 15.780 13.110 16.080 13.240 ;
        RECT 17.360 13.100 17.660 13.240 ;
        RECT 18.930 13.100 19.230 13.240 ;
        RECT 20.510 13.090 20.810 13.240 ;
        RECT 22.080 13.090 22.380 13.240 ;
        RECT 23.830 11.700 24.610 13.240 ;
        RECT 15.770 11.010 16.070 11.170 ;
        RECT 17.360 11.010 17.660 11.170 ;
        RECT 18.940 11.010 19.240 11.170 ;
        RECT 20.500 11.010 20.800 11.180 ;
        RECT 22.080 11.010 22.380 11.180 ;
        RECT 23.830 11.010 24.250 11.700 ;
        RECT 15.770 10.590 24.250 11.010 ;
        RECT 15.770 10.420 16.070 10.590 ;
        RECT 17.360 10.420 17.660 10.590 ;
        RECT 18.940 10.420 19.240 10.590 ;
        RECT 20.500 10.430 20.800 10.590 ;
        RECT 22.080 10.430 22.380 10.590 ;
      LAYER via2 ;
        RECT 16.850 106.390 17.390 106.930 ;
        RECT 5.015 78.505 5.505 78.995 ;
        RECT 10.725 78.455 11.215 78.945 ;
        RECT 16.850 34.670 17.390 35.210 ;
      LAYER met3 ;
        RECT 16.825 106.930 17.415 106.955 ;
        RECT 14.150 106.390 17.415 106.930 ;
        RECT 14.150 80.750 14.690 106.390 ;
        RECT 16.825 106.365 17.415 106.390 ;
        RECT 4.990 80.210 14.690 80.750 ;
        RECT 4.990 78.440 5.530 80.210 ;
        RECT 10.700 78.430 15.930 78.970 ;
        RECT 15.390 60.030 15.930 78.430 ;
        RECT 14.160 59.490 15.930 60.030 ;
        RECT 14.160 35.210 14.700 59.490 ;
        RECT 16.825 35.210 17.415 35.235 ;
        RECT 14.160 34.670 17.415 35.210 ;
        RECT 16.825 34.645 17.415 34.670 ;
  END
END audiodac_drv
END LIBRARY

