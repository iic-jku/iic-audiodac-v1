VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO audiodac
  CLASS BLOCK ;
  FOREIGN audiodac ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 2000.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END clk_i
  PIN ds_n_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 1996.000 750.170 2000.000 ;
    END
  END ds_n_o
  PIN ds_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 1996.000 250.150 2000.000 ;
    END
  END ds_o
  PIN fifo_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END fifo_ack_o
  PIN fifo_empty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END fifo_empty_o
  PIN fifo_full_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END fifo_full_o
  PIN fifo_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END fifo_i[0]
  PIN fifo_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END fifo_i[10]
  PIN fifo_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END fifo_i[11]
  PIN fifo_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END fifo_i[12]
  PIN fifo_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END fifo_i[13]
  PIN fifo_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END fifo_i[14]
  PIN fifo_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END fifo_i[15]
  PIN fifo_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END fifo_i[1]
  PIN fifo_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END fifo_i[2]
  PIN fifo_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END fifo_i[3]
  PIN fifo_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END fifo_i[4]
  PIN fifo_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END fifo_i[5]
  PIN fifo_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END fifo_i[6]
  PIN fifo_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END fifo_i[7]
  PIN fifo_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END fifo_i[8]
  PIN fifo_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END fifo_i[9]
  PIN fifo_rdy_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END fifo_rdy_i
  PIN mode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END mode_i
  PIN osr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END osr_i[0]
  PIN osr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END osr_i[1]
  PIN rst_n_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END rst_n_i
  PIN tst_fifo_loop_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END tst_fifo_loop_i
  PIN tst_sinegen_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 0.000 871.610 4.000 ;
    END
  END tst_sinegen_en_i
  PIN tst_sinegen_step_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END tst_sinegen_step_i[0]
  PIN tst_sinegen_step_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END tst_sinegen_step_i[1]
  PIN tst_sinegen_step_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.890 0.000 957.170 4.000 ;
    END
  END tst_sinegen_step_i[2]
  PIN tst_sinegen_step_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END tst_sinegen_step_i[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1988.560 ;
    END
  END vccd1
  PIN volume_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END volume_i[0]
  PIN volume_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END volume_i[1]
  PIN volume_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END volume_i[2]
  PIN volume_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END volume_i[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1988.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1988.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1986.905 994.250 1988.510 ;
        RECT 5.330 1981.465 994.250 1984.295 ;
        RECT 5.330 1976.025 994.250 1978.855 ;
        RECT 5.330 1970.585 994.250 1973.415 ;
        RECT 5.330 1965.145 994.250 1967.975 ;
        RECT 5.330 1959.705 994.250 1962.535 ;
        RECT 5.330 1954.265 994.250 1957.095 ;
        RECT 5.330 1948.825 994.250 1951.655 ;
        RECT 5.330 1943.385 994.250 1946.215 ;
        RECT 5.330 1937.945 994.250 1940.775 ;
        RECT 5.330 1932.505 994.250 1935.335 ;
        RECT 5.330 1927.065 994.250 1929.895 ;
        RECT 5.330 1921.625 994.250 1924.455 ;
        RECT 5.330 1916.185 994.250 1919.015 ;
        RECT 5.330 1910.745 994.250 1913.575 ;
        RECT 5.330 1905.305 994.250 1908.135 ;
        RECT 5.330 1899.865 994.250 1902.695 ;
        RECT 5.330 1894.425 994.250 1897.255 ;
        RECT 5.330 1888.985 994.250 1891.815 ;
        RECT 5.330 1883.545 994.250 1886.375 ;
        RECT 5.330 1878.105 994.250 1880.935 ;
        RECT 5.330 1872.665 994.250 1875.495 ;
        RECT 5.330 1867.225 994.250 1870.055 ;
        RECT 5.330 1861.785 994.250 1864.615 ;
        RECT 5.330 1856.345 994.250 1859.175 ;
        RECT 5.330 1850.905 994.250 1853.735 ;
        RECT 5.330 1845.465 994.250 1848.295 ;
        RECT 5.330 1840.025 994.250 1842.855 ;
        RECT 5.330 1834.585 994.250 1837.415 ;
        RECT 5.330 1829.145 994.250 1831.975 ;
        RECT 5.330 1823.705 994.250 1826.535 ;
        RECT 5.330 1818.265 994.250 1821.095 ;
        RECT 5.330 1812.825 994.250 1815.655 ;
        RECT 5.330 1807.385 994.250 1810.215 ;
        RECT 5.330 1801.945 994.250 1804.775 ;
        RECT 5.330 1796.505 994.250 1799.335 ;
        RECT 5.330 1791.065 994.250 1793.895 ;
        RECT 5.330 1785.625 994.250 1788.455 ;
        RECT 5.330 1780.185 994.250 1783.015 ;
        RECT 5.330 1774.745 994.250 1777.575 ;
        RECT 5.330 1769.305 994.250 1772.135 ;
        RECT 5.330 1763.865 994.250 1766.695 ;
        RECT 5.330 1758.425 994.250 1761.255 ;
        RECT 5.330 1752.985 994.250 1755.815 ;
        RECT 5.330 1747.545 994.250 1750.375 ;
        RECT 5.330 1742.105 994.250 1744.935 ;
        RECT 5.330 1736.665 994.250 1739.495 ;
        RECT 5.330 1731.225 994.250 1734.055 ;
        RECT 5.330 1725.785 994.250 1728.615 ;
        RECT 5.330 1720.345 994.250 1723.175 ;
        RECT 5.330 1714.905 994.250 1717.735 ;
        RECT 5.330 1709.465 994.250 1712.295 ;
        RECT 5.330 1704.025 994.250 1706.855 ;
        RECT 5.330 1698.585 994.250 1701.415 ;
        RECT 5.330 1693.145 994.250 1695.975 ;
        RECT 5.330 1687.705 994.250 1690.535 ;
        RECT 5.330 1682.265 994.250 1685.095 ;
        RECT 5.330 1676.825 994.250 1679.655 ;
        RECT 5.330 1671.385 994.250 1674.215 ;
        RECT 5.330 1665.945 994.250 1668.775 ;
        RECT 5.330 1660.505 994.250 1663.335 ;
        RECT 5.330 1655.065 994.250 1657.895 ;
        RECT 5.330 1649.625 994.250 1652.455 ;
        RECT 5.330 1644.185 994.250 1647.015 ;
        RECT 5.330 1638.745 994.250 1641.575 ;
        RECT 5.330 1633.305 994.250 1636.135 ;
        RECT 5.330 1627.865 994.250 1630.695 ;
        RECT 5.330 1622.425 994.250 1625.255 ;
        RECT 5.330 1616.985 994.250 1619.815 ;
        RECT 5.330 1611.545 994.250 1614.375 ;
        RECT 5.330 1606.105 994.250 1608.935 ;
        RECT 5.330 1600.665 994.250 1603.495 ;
        RECT 5.330 1595.225 994.250 1598.055 ;
        RECT 5.330 1589.785 994.250 1592.615 ;
        RECT 5.330 1584.345 994.250 1587.175 ;
        RECT 5.330 1578.905 994.250 1581.735 ;
        RECT 5.330 1573.465 994.250 1576.295 ;
        RECT 5.330 1568.025 994.250 1570.855 ;
        RECT 5.330 1562.585 994.250 1565.415 ;
        RECT 5.330 1557.145 994.250 1559.975 ;
        RECT 5.330 1551.705 994.250 1554.535 ;
        RECT 5.330 1546.265 994.250 1549.095 ;
        RECT 5.330 1540.825 994.250 1543.655 ;
        RECT 5.330 1535.385 994.250 1538.215 ;
        RECT 5.330 1529.945 994.250 1532.775 ;
        RECT 5.330 1524.505 994.250 1527.335 ;
        RECT 5.330 1519.065 994.250 1521.895 ;
        RECT 5.330 1513.625 994.250 1516.455 ;
        RECT 5.330 1508.185 994.250 1511.015 ;
        RECT 5.330 1502.745 994.250 1505.575 ;
        RECT 5.330 1497.305 994.250 1500.135 ;
        RECT 5.330 1491.865 994.250 1494.695 ;
        RECT 5.330 1486.425 994.250 1489.255 ;
        RECT 5.330 1480.985 994.250 1483.815 ;
        RECT 5.330 1475.545 994.250 1478.375 ;
        RECT 5.330 1470.105 994.250 1472.935 ;
        RECT 5.330 1464.665 994.250 1467.495 ;
        RECT 5.330 1459.225 994.250 1462.055 ;
        RECT 5.330 1453.785 994.250 1456.615 ;
        RECT 5.330 1448.345 994.250 1451.175 ;
        RECT 5.330 1442.905 994.250 1445.735 ;
        RECT 5.330 1437.465 994.250 1440.295 ;
        RECT 5.330 1432.025 994.250 1434.855 ;
        RECT 5.330 1426.585 994.250 1429.415 ;
        RECT 5.330 1421.145 994.250 1423.975 ;
        RECT 5.330 1415.705 994.250 1418.535 ;
        RECT 5.330 1410.265 994.250 1413.095 ;
        RECT 5.330 1404.825 994.250 1407.655 ;
        RECT 5.330 1399.385 994.250 1402.215 ;
        RECT 5.330 1393.945 994.250 1396.775 ;
        RECT 5.330 1388.505 994.250 1391.335 ;
        RECT 5.330 1383.065 994.250 1385.895 ;
        RECT 5.330 1377.625 994.250 1380.455 ;
        RECT 5.330 1372.185 994.250 1375.015 ;
        RECT 5.330 1366.745 994.250 1369.575 ;
        RECT 5.330 1361.305 994.250 1364.135 ;
        RECT 5.330 1355.865 994.250 1358.695 ;
        RECT 5.330 1350.425 994.250 1353.255 ;
        RECT 5.330 1344.985 994.250 1347.815 ;
        RECT 5.330 1339.545 994.250 1342.375 ;
        RECT 5.330 1334.105 994.250 1336.935 ;
        RECT 5.330 1328.665 994.250 1331.495 ;
        RECT 5.330 1323.225 994.250 1326.055 ;
        RECT 5.330 1317.785 994.250 1320.615 ;
        RECT 5.330 1312.345 994.250 1315.175 ;
        RECT 5.330 1306.905 994.250 1309.735 ;
        RECT 5.330 1301.465 994.250 1304.295 ;
        RECT 5.330 1296.025 994.250 1298.855 ;
        RECT 5.330 1290.585 994.250 1293.415 ;
        RECT 5.330 1285.145 994.250 1287.975 ;
        RECT 5.330 1279.705 994.250 1282.535 ;
        RECT 5.330 1274.265 994.250 1277.095 ;
        RECT 5.330 1268.825 994.250 1271.655 ;
        RECT 5.330 1263.385 994.250 1266.215 ;
        RECT 5.330 1257.945 994.250 1260.775 ;
        RECT 5.330 1252.505 994.250 1255.335 ;
        RECT 5.330 1247.065 994.250 1249.895 ;
        RECT 5.330 1241.625 994.250 1244.455 ;
        RECT 5.330 1236.185 994.250 1239.015 ;
        RECT 5.330 1230.745 994.250 1233.575 ;
        RECT 5.330 1225.305 994.250 1228.135 ;
        RECT 5.330 1219.865 994.250 1222.695 ;
        RECT 5.330 1214.425 994.250 1217.255 ;
        RECT 5.330 1208.985 994.250 1211.815 ;
        RECT 5.330 1203.545 994.250 1206.375 ;
        RECT 5.330 1198.105 994.250 1200.935 ;
        RECT 5.330 1192.665 994.250 1195.495 ;
        RECT 5.330 1187.225 994.250 1190.055 ;
        RECT 5.330 1181.785 994.250 1184.615 ;
        RECT 5.330 1176.345 994.250 1179.175 ;
        RECT 5.330 1170.905 994.250 1173.735 ;
        RECT 5.330 1165.465 994.250 1168.295 ;
        RECT 5.330 1160.025 994.250 1162.855 ;
        RECT 5.330 1154.585 994.250 1157.415 ;
        RECT 5.330 1149.145 994.250 1151.975 ;
        RECT 5.330 1143.705 994.250 1146.535 ;
        RECT 5.330 1138.265 994.250 1141.095 ;
        RECT 5.330 1132.825 994.250 1135.655 ;
        RECT 5.330 1127.385 994.250 1130.215 ;
        RECT 5.330 1121.945 994.250 1124.775 ;
        RECT 5.330 1116.505 994.250 1119.335 ;
        RECT 5.330 1111.065 994.250 1113.895 ;
        RECT 5.330 1105.625 994.250 1108.455 ;
        RECT 5.330 1100.185 994.250 1103.015 ;
        RECT 5.330 1094.745 994.250 1097.575 ;
        RECT 5.330 1089.305 994.250 1092.135 ;
        RECT 5.330 1083.865 994.250 1086.695 ;
        RECT 5.330 1078.425 994.250 1081.255 ;
        RECT 5.330 1072.985 994.250 1075.815 ;
        RECT 5.330 1067.545 994.250 1070.375 ;
        RECT 5.330 1062.105 994.250 1064.935 ;
        RECT 5.330 1056.665 994.250 1059.495 ;
        RECT 5.330 1051.225 994.250 1054.055 ;
        RECT 5.330 1045.785 994.250 1048.615 ;
        RECT 5.330 1040.345 994.250 1043.175 ;
        RECT 5.330 1034.905 994.250 1037.735 ;
        RECT 5.330 1029.465 994.250 1032.295 ;
        RECT 5.330 1024.025 994.250 1026.855 ;
        RECT 5.330 1018.585 994.250 1021.415 ;
        RECT 5.330 1013.145 994.250 1015.975 ;
        RECT 5.330 1007.705 994.250 1010.535 ;
        RECT 5.330 1002.265 994.250 1005.095 ;
        RECT 5.330 996.825 994.250 999.655 ;
        RECT 5.330 991.385 994.250 994.215 ;
        RECT 5.330 985.945 994.250 988.775 ;
        RECT 5.330 980.505 994.250 983.335 ;
        RECT 5.330 975.065 994.250 977.895 ;
        RECT 5.330 969.625 994.250 972.455 ;
        RECT 5.330 964.185 994.250 967.015 ;
        RECT 5.330 958.745 994.250 961.575 ;
        RECT 5.330 953.305 994.250 956.135 ;
        RECT 5.330 947.865 994.250 950.695 ;
        RECT 5.330 942.425 994.250 945.255 ;
        RECT 5.330 936.985 994.250 939.815 ;
        RECT 5.330 931.545 994.250 934.375 ;
        RECT 5.330 926.105 994.250 928.935 ;
        RECT 5.330 920.665 994.250 923.495 ;
        RECT 5.330 915.225 994.250 918.055 ;
        RECT 5.330 909.785 994.250 912.615 ;
        RECT 5.330 904.345 994.250 907.175 ;
        RECT 5.330 898.905 994.250 901.735 ;
        RECT 5.330 893.465 994.250 896.295 ;
        RECT 5.330 888.025 994.250 890.855 ;
        RECT 5.330 882.585 994.250 885.415 ;
        RECT 5.330 877.145 994.250 879.975 ;
        RECT 5.330 871.705 994.250 874.535 ;
        RECT 5.330 866.265 994.250 869.095 ;
        RECT 5.330 860.825 994.250 863.655 ;
        RECT 5.330 855.385 994.250 858.215 ;
        RECT 5.330 849.945 994.250 852.775 ;
        RECT 5.330 844.505 994.250 847.335 ;
        RECT 5.330 839.065 994.250 841.895 ;
        RECT 5.330 833.625 994.250 836.455 ;
        RECT 5.330 828.185 994.250 831.015 ;
        RECT 5.330 822.745 994.250 825.575 ;
        RECT 5.330 817.305 994.250 820.135 ;
        RECT 5.330 811.865 994.250 814.695 ;
        RECT 5.330 806.425 994.250 809.255 ;
        RECT 5.330 800.985 994.250 803.815 ;
        RECT 5.330 795.545 994.250 798.375 ;
        RECT 5.330 790.105 994.250 792.935 ;
        RECT 5.330 784.665 994.250 787.495 ;
        RECT 5.330 779.225 994.250 782.055 ;
        RECT 5.330 773.785 994.250 776.615 ;
        RECT 5.330 768.345 994.250 771.175 ;
        RECT 5.330 762.905 994.250 765.735 ;
        RECT 5.330 757.465 994.250 760.295 ;
        RECT 5.330 752.025 994.250 754.855 ;
        RECT 5.330 746.585 994.250 749.415 ;
        RECT 5.330 741.145 994.250 743.975 ;
        RECT 5.330 735.705 994.250 738.535 ;
        RECT 5.330 730.265 994.250 733.095 ;
        RECT 5.330 724.825 994.250 727.655 ;
        RECT 5.330 719.385 994.250 722.215 ;
        RECT 5.330 713.945 994.250 716.775 ;
        RECT 5.330 708.505 994.250 711.335 ;
        RECT 5.330 703.065 994.250 705.895 ;
        RECT 5.330 697.625 994.250 700.455 ;
        RECT 5.330 692.185 994.250 695.015 ;
        RECT 5.330 686.745 994.250 689.575 ;
        RECT 5.330 681.305 994.250 684.135 ;
        RECT 5.330 675.865 994.250 678.695 ;
        RECT 5.330 670.425 994.250 673.255 ;
        RECT 5.330 664.985 994.250 667.815 ;
        RECT 5.330 659.545 994.250 662.375 ;
        RECT 5.330 654.105 994.250 656.935 ;
        RECT 5.330 648.665 994.250 651.495 ;
        RECT 5.330 643.225 994.250 646.055 ;
        RECT 5.330 637.785 994.250 640.615 ;
        RECT 5.330 632.345 994.250 635.175 ;
        RECT 5.330 626.905 994.250 629.735 ;
        RECT 5.330 621.465 994.250 624.295 ;
        RECT 5.330 616.025 994.250 618.855 ;
        RECT 5.330 610.585 994.250 613.415 ;
        RECT 5.330 605.145 994.250 607.975 ;
        RECT 5.330 599.705 994.250 602.535 ;
        RECT 5.330 594.265 994.250 597.095 ;
        RECT 5.330 588.825 994.250 591.655 ;
        RECT 5.330 583.385 994.250 586.215 ;
        RECT 5.330 577.945 994.250 580.775 ;
        RECT 5.330 572.505 994.250 575.335 ;
        RECT 5.330 567.065 994.250 569.895 ;
        RECT 5.330 561.625 994.250 564.455 ;
        RECT 5.330 556.185 994.250 559.015 ;
        RECT 5.330 550.745 994.250 553.575 ;
        RECT 5.330 545.305 994.250 548.135 ;
        RECT 5.330 539.865 994.250 542.695 ;
        RECT 5.330 534.425 994.250 537.255 ;
        RECT 5.330 528.985 994.250 531.815 ;
        RECT 5.330 523.545 994.250 526.375 ;
        RECT 5.330 518.105 994.250 520.935 ;
        RECT 5.330 512.665 994.250 515.495 ;
        RECT 5.330 507.225 994.250 510.055 ;
        RECT 5.330 501.785 994.250 504.615 ;
        RECT 5.330 496.345 994.250 499.175 ;
        RECT 5.330 490.905 994.250 493.735 ;
        RECT 5.330 485.465 994.250 488.295 ;
        RECT 5.330 480.025 994.250 482.855 ;
        RECT 5.330 474.585 994.250 477.415 ;
        RECT 5.330 469.145 994.250 471.975 ;
        RECT 5.330 463.705 994.250 466.535 ;
        RECT 5.330 458.265 994.250 461.095 ;
        RECT 5.330 452.825 994.250 455.655 ;
        RECT 5.330 447.385 994.250 450.215 ;
        RECT 5.330 441.945 994.250 444.775 ;
        RECT 5.330 436.505 994.250 439.335 ;
        RECT 5.330 431.065 994.250 433.895 ;
        RECT 5.330 425.625 994.250 428.455 ;
        RECT 5.330 420.185 994.250 423.015 ;
        RECT 5.330 414.745 994.250 417.575 ;
        RECT 5.330 409.305 994.250 412.135 ;
        RECT 5.330 403.865 994.250 406.695 ;
        RECT 5.330 398.425 994.250 401.255 ;
        RECT 5.330 392.985 994.250 395.815 ;
        RECT 5.330 387.545 994.250 390.375 ;
        RECT 5.330 382.105 994.250 384.935 ;
        RECT 5.330 376.665 994.250 379.495 ;
        RECT 5.330 371.225 994.250 374.055 ;
        RECT 5.330 365.785 994.250 368.615 ;
        RECT 5.330 360.345 994.250 363.175 ;
        RECT 5.330 354.905 994.250 357.735 ;
        RECT 5.330 349.465 994.250 352.295 ;
        RECT 5.330 344.025 994.250 346.855 ;
        RECT 5.330 338.585 994.250 341.415 ;
        RECT 5.330 333.145 994.250 335.975 ;
        RECT 5.330 327.705 994.250 330.535 ;
        RECT 5.330 322.265 994.250 325.095 ;
        RECT 5.330 316.825 994.250 319.655 ;
        RECT 5.330 311.385 994.250 314.215 ;
        RECT 5.330 305.945 994.250 308.775 ;
        RECT 5.330 300.505 994.250 303.335 ;
        RECT 5.330 295.065 994.250 297.895 ;
        RECT 5.330 289.625 994.250 292.455 ;
        RECT 5.330 284.185 994.250 287.015 ;
        RECT 5.330 278.745 994.250 281.575 ;
        RECT 5.330 273.305 994.250 276.135 ;
        RECT 5.330 267.865 994.250 270.695 ;
        RECT 5.330 262.425 994.250 265.255 ;
        RECT 5.330 256.985 994.250 259.815 ;
        RECT 5.330 251.545 994.250 254.375 ;
        RECT 5.330 246.105 994.250 248.935 ;
        RECT 5.330 240.665 994.250 243.495 ;
        RECT 5.330 235.225 994.250 238.055 ;
        RECT 5.330 229.785 994.250 232.615 ;
        RECT 5.330 224.345 994.250 227.175 ;
        RECT 5.330 218.905 994.250 221.735 ;
        RECT 5.330 213.465 994.250 216.295 ;
        RECT 5.330 208.025 994.250 210.855 ;
        RECT 5.330 202.585 994.250 205.415 ;
        RECT 5.330 197.145 994.250 199.975 ;
        RECT 5.330 191.705 994.250 194.535 ;
        RECT 5.330 186.265 994.250 189.095 ;
        RECT 5.330 180.825 994.250 183.655 ;
        RECT 5.330 175.385 994.250 178.215 ;
        RECT 5.330 169.945 994.250 172.775 ;
        RECT 5.330 164.505 994.250 167.335 ;
        RECT 5.330 159.065 994.250 161.895 ;
        RECT 5.330 153.625 994.250 156.455 ;
        RECT 5.330 148.185 994.250 151.015 ;
        RECT 5.330 142.745 994.250 145.575 ;
        RECT 5.330 137.305 994.250 140.135 ;
        RECT 5.330 131.865 994.250 134.695 ;
        RECT 5.330 126.425 994.250 129.255 ;
        RECT 5.330 120.985 994.250 123.815 ;
        RECT 5.330 115.545 994.250 118.375 ;
        RECT 5.330 110.105 994.250 112.935 ;
        RECT 5.330 104.665 994.250 107.495 ;
        RECT 5.330 99.225 994.250 102.055 ;
        RECT 5.330 93.785 994.250 96.615 ;
        RECT 5.330 88.345 994.250 91.175 ;
        RECT 5.330 82.905 994.250 85.735 ;
        RECT 5.330 77.465 994.250 80.295 ;
        RECT 5.330 72.025 994.250 74.855 ;
        RECT 5.330 66.585 994.250 69.415 ;
        RECT 5.330 61.145 994.250 63.975 ;
        RECT 5.330 55.705 994.250 58.535 ;
        RECT 5.330 50.265 994.250 53.095 ;
        RECT 5.330 44.825 994.250 47.655 ;
        RECT 5.330 39.385 994.250 42.215 ;
        RECT 5.330 33.945 994.250 36.775 ;
        RECT 5.330 28.505 994.250 31.335 ;
        RECT 5.330 23.065 994.250 25.895 ;
        RECT 5.330 17.625 994.250 20.455 ;
        RECT 5.330 12.185 994.250 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 994.060 1988.405 ;
      LAYER met1 ;
        RECT 5.520 10.240 994.060 1988.560 ;
      LAYER met2 ;
        RECT 14.360 1995.720 249.590 1996.000 ;
        RECT 250.430 1995.720 749.610 1996.000 ;
        RECT 750.450 1995.720 989.820 1996.000 ;
        RECT 14.360 4.280 989.820 1995.720 ;
        RECT 14.910 3.670 42.590 4.280 ;
        RECT 43.430 3.670 71.110 4.280 ;
        RECT 71.950 3.670 99.630 4.280 ;
        RECT 100.470 3.670 128.150 4.280 ;
        RECT 128.990 3.670 156.670 4.280 ;
        RECT 157.510 3.670 185.190 4.280 ;
        RECT 186.030 3.670 213.710 4.280 ;
        RECT 214.550 3.670 242.230 4.280 ;
        RECT 243.070 3.670 271.210 4.280 ;
        RECT 272.050 3.670 299.730 4.280 ;
        RECT 300.570 3.670 328.250 4.280 ;
        RECT 329.090 3.670 356.770 4.280 ;
        RECT 357.610 3.670 385.290 4.280 ;
        RECT 386.130 3.670 413.810 4.280 ;
        RECT 414.650 3.670 442.330 4.280 ;
        RECT 443.170 3.670 470.850 4.280 ;
        RECT 471.690 3.670 499.370 4.280 ;
        RECT 500.210 3.670 528.350 4.280 ;
        RECT 529.190 3.670 556.870 4.280 ;
        RECT 557.710 3.670 585.390 4.280 ;
        RECT 586.230 3.670 613.910 4.280 ;
        RECT 614.750 3.670 642.430 4.280 ;
        RECT 643.270 3.670 670.950 4.280 ;
        RECT 671.790 3.670 699.470 4.280 ;
        RECT 700.310 3.670 727.990 4.280 ;
        RECT 728.830 3.670 756.510 4.280 ;
        RECT 757.350 3.670 785.490 4.280 ;
        RECT 786.330 3.670 814.010 4.280 ;
        RECT 814.850 3.670 842.530 4.280 ;
        RECT 843.370 3.670 871.050 4.280 ;
        RECT 871.890 3.670 899.570 4.280 ;
        RECT 900.410 3.670 928.090 4.280 ;
        RECT 928.930 3.670 956.610 4.280 ;
        RECT 957.450 3.670 985.130 4.280 ;
        RECT 985.970 3.670 989.820 4.280 ;
      LAYER met3 ;
        RECT 21.040 10.715 944.240 1988.485 ;
      LAYER met4 ;
        RECT 171.415 17.175 174.240 1970.465 ;
        RECT 176.640 17.175 251.040 1970.465 ;
        RECT 253.440 17.175 327.840 1970.465 ;
        RECT 330.240 17.175 404.640 1970.465 ;
        RECT 407.040 17.175 481.440 1970.465 ;
        RECT 483.840 17.175 558.240 1970.465 ;
        RECT 560.640 17.175 635.040 1970.465 ;
        RECT 637.440 17.175 711.840 1970.465 ;
        RECT 714.240 17.175 788.640 1970.465 ;
        RECT 791.040 17.175 865.440 1970.465 ;
        RECT 867.840 17.175 868.185 1970.465 ;
  END
END audiodac
END LIBRARY

