magic
tech sky130A
magscale 1 2
timestamp 1644774117
<< obsli1 >>
rect 1104 2159 398820 397681
<< obsm1 >>
rect 1104 1640 398820 397712
<< metal2 >>
rect 1582 399200 1638 400000
rect 4802 399200 4858 400000
rect 8022 399200 8078 400000
rect 11334 399200 11390 400000
rect 14554 399200 14610 400000
rect 17774 399200 17830 400000
rect 21086 399200 21142 400000
rect 24306 399200 24362 400000
rect 27526 399200 27582 400000
rect 30838 399200 30894 400000
rect 34058 399200 34114 400000
rect 37278 399200 37334 400000
rect 40590 399200 40646 400000
rect 43810 399200 43866 400000
rect 47030 399200 47086 400000
rect 50342 399200 50398 400000
rect 53562 399200 53618 400000
rect 56782 399200 56838 400000
rect 60094 399200 60150 400000
rect 63314 399200 63370 400000
rect 66534 399200 66590 400000
rect 69846 399200 69902 400000
rect 73066 399200 73122 400000
rect 76378 399200 76434 400000
rect 79598 399200 79654 400000
rect 82818 399200 82874 400000
rect 86130 399200 86186 400000
rect 89350 399200 89406 400000
rect 92570 399200 92626 400000
rect 95882 399200 95938 400000
rect 99102 399200 99158 400000
rect 102322 399200 102378 400000
rect 105634 399200 105690 400000
rect 108854 399200 108910 400000
rect 112074 399200 112130 400000
rect 115386 399200 115442 400000
rect 118606 399200 118662 400000
rect 121826 399200 121882 400000
rect 125138 399200 125194 400000
rect 128358 399200 128414 400000
rect 131578 399200 131634 400000
rect 134890 399200 134946 400000
rect 138110 399200 138166 400000
rect 141422 399200 141478 400000
rect 144642 399200 144698 400000
rect 147862 399200 147918 400000
rect 151174 399200 151230 400000
rect 154394 399200 154450 400000
rect 157614 399200 157670 400000
rect 160926 399200 160982 400000
rect 164146 399200 164202 400000
rect 167366 399200 167422 400000
rect 170678 399200 170734 400000
rect 173898 399200 173954 400000
rect 177118 399200 177174 400000
rect 180430 399200 180486 400000
rect 183650 399200 183706 400000
rect 186870 399200 186926 400000
rect 190182 399200 190238 400000
rect 193402 399200 193458 400000
rect 196622 399200 196678 400000
rect 199934 399200 199990 400000
rect 203154 399200 203210 400000
rect 206466 399200 206522 400000
rect 209686 399200 209742 400000
rect 212906 399200 212962 400000
rect 216218 399200 216274 400000
rect 219438 399200 219494 400000
rect 222658 399200 222714 400000
rect 225970 399200 226026 400000
rect 229190 399200 229246 400000
rect 232410 399200 232466 400000
rect 235722 399200 235778 400000
rect 238942 399200 238998 400000
rect 242162 399200 242218 400000
rect 245474 399200 245530 400000
rect 248694 399200 248750 400000
rect 251914 399200 251970 400000
rect 255226 399200 255282 400000
rect 258446 399200 258502 400000
rect 261666 399200 261722 400000
rect 264978 399200 265034 400000
rect 268198 399200 268254 400000
rect 271510 399200 271566 400000
rect 274730 399200 274786 400000
rect 277950 399200 278006 400000
rect 281262 399200 281318 400000
rect 284482 399200 284538 400000
rect 287702 399200 287758 400000
rect 291014 399200 291070 400000
rect 294234 399200 294290 400000
rect 297454 399200 297510 400000
rect 300766 399200 300822 400000
rect 303986 399200 304042 400000
rect 307206 399200 307262 400000
rect 310518 399200 310574 400000
rect 313738 399200 313794 400000
rect 316958 399200 317014 400000
rect 320270 399200 320326 400000
rect 323490 399200 323546 400000
rect 326710 399200 326766 400000
rect 330022 399200 330078 400000
rect 333242 399200 333298 400000
rect 336554 399200 336610 400000
rect 339774 399200 339830 400000
rect 342994 399200 343050 400000
rect 346306 399200 346362 400000
rect 349526 399200 349582 400000
rect 352746 399200 352802 400000
rect 356058 399200 356114 400000
rect 359278 399200 359334 400000
rect 362498 399200 362554 400000
rect 365810 399200 365866 400000
rect 369030 399200 369086 400000
rect 372250 399200 372306 400000
rect 375562 399200 375618 400000
rect 378782 399200 378838 400000
rect 382002 399200 382058 400000
rect 385314 399200 385370 400000
rect 388534 399200 388590 400000
rect 391754 399200 391810 400000
rect 395066 399200 395122 400000
rect 398286 399200 398342 400000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2686 0 2742 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 5078 0 5134 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7470 0 7526 800
rect 8206 0 8262 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10598 0 10654 800
rect 11426 0 11482 800
rect 12162 0 12218 800
rect 12990 0 13046 800
rect 13726 0 13782 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18510 0 18566 800
rect 19246 0 19302 800
rect 20074 0 20130 800
rect 20810 0 20866 800
rect 21638 0 21694 800
rect 22466 0 22522 800
rect 23202 0 23258 800
rect 24030 0 24086 800
rect 24766 0 24822 800
rect 25594 0 25650 800
rect 26422 0 26478 800
rect 27158 0 27214 800
rect 27986 0 28042 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30286 0 30342 800
rect 31114 0 31170 800
rect 31942 0 31998 800
rect 32678 0 32734 800
rect 33506 0 33562 800
rect 34242 0 34298 800
rect 35070 0 35126 800
rect 35806 0 35862 800
rect 36634 0 36690 800
rect 37462 0 37518 800
rect 38198 0 38254 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40590 0 40646 800
rect 41326 0 41382 800
rect 42154 0 42210 800
rect 42982 0 43038 800
rect 43718 0 43774 800
rect 44546 0 44602 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46846 0 46902 800
rect 47674 0 47730 800
rect 48502 0 48558 800
rect 49238 0 49294 800
rect 50066 0 50122 800
rect 50802 0 50858 800
rect 51630 0 51686 800
rect 52458 0 52514 800
rect 53194 0 53250 800
rect 54022 0 54078 800
rect 54758 0 54814 800
rect 55586 0 55642 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60278 0 60334 800
rect 61106 0 61162 800
rect 61842 0 61898 800
rect 62670 0 62726 800
rect 63498 0 63554 800
rect 64234 0 64290 800
rect 65062 0 65118 800
rect 65798 0 65854 800
rect 66626 0 66682 800
rect 67362 0 67418 800
rect 68190 0 68246 800
rect 69018 0 69074 800
rect 69754 0 69810 800
rect 70582 0 70638 800
rect 71318 0 71374 800
rect 72146 0 72202 800
rect 72882 0 72938 800
rect 73710 0 73766 800
rect 74538 0 74594 800
rect 75274 0 75330 800
rect 76102 0 76158 800
rect 76838 0 76894 800
rect 77666 0 77722 800
rect 78494 0 78550 800
rect 79230 0 79286 800
rect 80058 0 80114 800
rect 80794 0 80850 800
rect 81622 0 81678 800
rect 82358 0 82414 800
rect 83186 0 83242 800
rect 84014 0 84070 800
rect 84750 0 84806 800
rect 85578 0 85634 800
rect 86314 0 86370 800
rect 87142 0 87198 800
rect 87878 0 87934 800
rect 88706 0 88762 800
rect 89534 0 89590 800
rect 90270 0 90326 800
rect 91098 0 91154 800
rect 91834 0 91890 800
rect 92662 0 92718 800
rect 93398 0 93454 800
rect 94226 0 94282 800
rect 95054 0 95110 800
rect 95790 0 95846 800
rect 96618 0 96674 800
rect 97354 0 97410 800
rect 98182 0 98238 800
rect 98918 0 98974 800
rect 99746 0 99802 800
rect 100574 0 100630 800
rect 101310 0 101366 800
rect 102138 0 102194 800
rect 102874 0 102930 800
rect 103702 0 103758 800
rect 104530 0 104586 800
rect 105266 0 105322 800
rect 106094 0 106150 800
rect 106830 0 106886 800
rect 107658 0 107714 800
rect 108394 0 108450 800
rect 109222 0 109278 800
rect 110050 0 110106 800
rect 110786 0 110842 800
rect 111614 0 111670 800
rect 112350 0 112406 800
rect 113178 0 113234 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115570 0 115626 800
rect 116306 0 116362 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118698 0 118754 800
rect 119434 0 119490 800
rect 120262 0 120318 800
rect 121090 0 121146 800
rect 121826 0 121882 800
rect 122654 0 122710 800
rect 123390 0 123446 800
rect 124218 0 124274 800
rect 124954 0 125010 800
rect 125782 0 125838 800
rect 126610 0 126666 800
rect 127346 0 127402 800
rect 128174 0 128230 800
rect 128910 0 128966 800
rect 129738 0 129794 800
rect 130566 0 130622 800
rect 131302 0 131358 800
rect 132130 0 132186 800
rect 132866 0 132922 800
rect 133694 0 133750 800
rect 134430 0 134486 800
rect 135258 0 135314 800
rect 136086 0 136142 800
rect 136822 0 136878 800
rect 137650 0 137706 800
rect 138386 0 138442 800
rect 139214 0 139270 800
rect 139950 0 140006 800
rect 140778 0 140834 800
rect 141606 0 141662 800
rect 142342 0 142398 800
rect 143170 0 143226 800
rect 143906 0 143962 800
rect 144734 0 144790 800
rect 145470 0 145526 800
rect 146298 0 146354 800
rect 147126 0 147182 800
rect 147862 0 147918 800
rect 148690 0 148746 800
rect 149426 0 149482 800
rect 150254 0 150310 800
rect 151082 0 151138 800
rect 151818 0 151874 800
rect 152646 0 152702 800
rect 153382 0 153438 800
rect 154210 0 154266 800
rect 154946 0 155002 800
rect 155774 0 155830 800
rect 156602 0 156658 800
rect 157338 0 157394 800
rect 158166 0 158222 800
rect 158902 0 158958 800
rect 159730 0 159786 800
rect 160466 0 160522 800
rect 161294 0 161350 800
rect 162122 0 162178 800
rect 162858 0 162914 800
rect 163686 0 163742 800
rect 164422 0 164478 800
rect 165250 0 165306 800
rect 165986 0 166042 800
rect 166814 0 166870 800
rect 167642 0 167698 800
rect 168378 0 168434 800
rect 169206 0 169262 800
rect 169942 0 169998 800
rect 170770 0 170826 800
rect 171506 0 171562 800
rect 172334 0 172390 800
rect 173162 0 173218 800
rect 173898 0 173954 800
rect 174726 0 174782 800
rect 175462 0 175518 800
rect 176290 0 176346 800
rect 177118 0 177174 800
rect 177854 0 177910 800
rect 178682 0 178738 800
rect 179418 0 179474 800
rect 180246 0 180302 800
rect 180982 0 181038 800
rect 181810 0 181866 800
rect 182638 0 182694 800
rect 183374 0 183430 800
rect 184202 0 184258 800
rect 184938 0 184994 800
rect 185766 0 185822 800
rect 186502 0 186558 800
rect 187330 0 187386 800
rect 188158 0 188214 800
rect 188894 0 188950 800
rect 189722 0 189778 800
rect 190458 0 190514 800
rect 191286 0 191342 800
rect 192022 0 192078 800
rect 192850 0 192906 800
rect 193678 0 193734 800
rect 194414 0 194470 800
rect 195242 0 195298 800
rect 195978 0 196034 800
rect 196806 0 196862 800
rect 197542 0 197598 800
rect 198370 0 198426 800
rect 199198 0 199254 800
rect 199934 0 199990 800
rect 200762 0 200818 800
rect 201498 0 201554 800
rect 202326 0 202382 800
rect 203154 0 203210 800
rect 203890 0 203946 800
rect 204718 0 204774 800
rect 205454 0 205510 800
rect 206282 0 206338 800
rect 207018 0 207074 800
rect 207846 0 207902 800
rect 208674 0 208730 800
rect 209410 0 209466 800
rect 210238 0 210294 800
rect 210974 0 211030 800
rect 211802 0 211858 800
rect 212538 0 212594 800
rect 213366 0 213422 800
rect 214194 0 214250 800
rect 214930 0 214986 800
rect 215758 0 215814 800
rect 216494 0 216550 800
rect 217322 0 217378 800
rect 218058 0 218114 800
rect 218886 0 218942 800
rect 219714 0 219770 800
rect 220450 0 220506 800
rect 221278 0 221334 800
rect 222014 0 222070 800
rect 222842 0 222898 800
rect 223578 0 223634 800
rect 224406 0 224462 800
rect 225234 0 225290 800
rect 225970 0 226026 800
rect 226798 0 226854 800
rect 227534 0 227590 800
rect 228362 0 228418 800
rect 229190 0 229246 800
rect 229926 0 229982 800
rect 230754 0 230810 800
rect 231490 0 231546 800
rect 232318 0 232374 800
rect 233054 0 233110 800
rect 233882 0 233938 800
rect 234710 0 234766 800
rect 235446 0 235502 800
rect 236274 0 236330 800
rect 237010 0 237066 800
rect 237838 0 237894 800
rect 238574 0 238630 800
rect 239402 0 239458 800
rect 240230 0 240286 800
rect 240966 0 241022 800
rect 241794 0 241850 800
rect 242530 0 242586 800
rect 243358 0 243414 800
rect 244094 0 244150 800
rect 244922 0 244978 800
rect 245750 0 245806 800
rect 246486 0 246542 800
rect 247314 0 247370 800
rect 248050 0 248106 800
rect 248878 0 248934 800
rect 249614 0 249670 800
rect 250442 0 250498 800
rect 251270 0 251326 800
rect 252006 0 252062 800
rect 252834 0 252890 800
rect 253570 0 253626 800
rect 254398 0 254454 800
rect 255226 0 255282 800
rect 255962 0 256018 800
rect 256790 0 256846 800
rect 257526 0 257582 800
rect 258354 0 258410 800
rect 259090 0 259146 800
rect 259918 0 259974 800
rect 260746 0 260802 800
rect 261482 0 261538 800
rect 262310 0 262366 800
rect 263046 0 263102 800
rect 263874 0 263930 800
rect 264610 0 264666 800
rect 265438 0 265494 800
rect 266266 0 266322 800
rect 267002 0 267058 800
rect 267830 0 267886 800
rect 268566 0 268622 800
rect 269394 0 269450 800
rect 270130 0 270186 800
rect 270958 0 271014 800
rect 271786 0 271842 800
rect 272522 0 272578 800
rect 273350 0 273406 800
rect 274086 0 274142 800
rect 274914 0 274970 800
rect 275742 0 275798 800
rect 276478 0 276534 800
rect 277306 0 277362 800
rect 278042 0 278098 800
rect 278870 0 278926 800
rect 279606 0 279662 800
rect 280434 0 280490 800
rect 281262 0 281318 800
rect 281998 0 282054 800
rect 282826 0 282882 800
rect 283562 0 283618 800
rect 284390 0 284446 800
rect 285126 0 285182 800
rect 285954 0 286010 800
rect 286782 0 286838 800
rect 287518 0 287574 800
rect 288346 0 288402 800
rect 289082 0 289138 800
rect 289910 0 289966 800
rect 290646 0 290702 800
rect 291474 0 291530 800
rect 292302 0 292358 800
rect 293038 0 293094 800
rect 293866 0 293922 800
rect 294602 0 294658 800
rect 295430 0 295486 800
rect 296166 0 296222 800
rect 296994 0 297050 800
rect 297822 0 297878 800
rect 298558 0 298614 800
rect 299386 0 299442 800
rect 300122 0 300178 800
rect 300950 0 301006 800
rect 301778 0 301834 800
rect 302514 0 302570 800
rect 303342 0 303398 800
rect 304078 0 304134 800
rect 304906 0 304962 800
rect 305642 0 305698 800
rect 306470 0 306526 800
rect 307298 0 307354 800
rect 308034 0 308090 800
rect 308862 0 308918 800
rect 309598 0 309654 800
rect 310426 0 310482 800
rect 311162 0 311218 800
rect 311990 0 312046 800
rect 312818 0 312874 800
rect 313554 0 313610 800
rect 314382 0 314438 800
rect 315118 0 315174 800
rect 315946 0 316002 800
rect 316682 0 316738 800
rect 317510 0 317566 800
rect 318338 0 318394 800
rect 319074 0 319130 800
rect 319902 0 319958 800
rect 320638 0 320694 800
rect 321466 0 321522 800
rect 322202 0 322258 800
rect 323030 0 323086 800
rect 323858 0 323914 800
rect 324594 0 324650 800
rect 325422 0 325478 800
rect 326158 0 326214 800
rect 326986 0 327042 800
rect 327814 0 327870 800
rect 328550 0 328606 800
rect 329378 0 329434 800
rect 330114 0 330170 800
rect 330942 0 330998 800
rect 331678 0 331734 800
rect 332506 0 332562 800
rect 333334 0 333390 800
rect 334070 0 334126 800
rect 334898 0 334954 800
rect 335634 0 335690 800
rect 336462 0 336518 800
rect 337198 0 337254 800
rect 338026 0 338082 800
rect 338854 0 338910 800
rect 339590 0 339646 800
rect 340418 0 340474 800
rect 341154 0 341210 800
rect 341982 0 342038 800
rect 342718 0 342774 800
rect 343546 0 343602 800
rect 344374 0 344430 800
rect 345110 0 345166 800
rect 345938 0 345994 800
rect 346674 0 346730 800
rect 347502 0 347558 800
rect 348238 0 348294 800
rect 349066 0 349122 800
rect 349894 0 349950 800
rect 350630 0 350686 800
rect 351458 0 351514 800
rect 352194 0 352250 800
rect 353022 0 353078 800
rect 353850 0 353906 800
rect 354586 0 354642 800
rect 355414 0 355470 800
rect 356150 0 356206 800
rect 356978 0 357034 800
rect 357714 0 357770 800
rect 358542 0 358598 800
rect 359370 0 359426 800
rect 360106 0 360162 800
rect 360934 0 360990 800
rect 361670 0 361726 800
rect 362498 0 362554 800
rect 363234 0 363290 800
rect 364062 0 364118 800
rect 364890 0 364946 800
rect 365626 0 365682 800
rect 366454 0 366510 800
rect 367190 0 367246 800
rect 368018 0 368074 800
rect 368754 0 368810 800
rect 369582 0 369638 800
rect 370410 0 370466 800
rect 371146 0 371202 800
rect 371974 0 372030 800
rect 372710 0 372766 800
rect 373538 0 373594 800
rect 374274 0 374330 800
rect 375102 0 375158 800
rect 375930 0 375986 800
rect 376666 0 376722 800
rect 377494 0 377550 800
rect 378230 0 378286 800
rect 379058 0 379114 800
rect 379886 0 379942 800
rect 380622 0 380678 800
rect 381450 0 381506 800
rect 382186 0 382242 800
rect 383014 0 383070 800
rect 383750 0 383806 800
rect 384578 0 384634 800
rect 385406 0 385462 800
rect 386142 0 386198 800
rect 386970 0 387026 800
rect 387706 0 387762 800
rect 388534 0 388590 800
rect 389270 0 389326 800
rect 390098 0 390154 800
rect 390926 0 390982 800
rect 391662 0 391718 800
rect 392490 0 392546 800
rect 393226 0 393282 800
rect 394054 0 394110 800
rect 394790 0 394846 800
rect 395618 0 395674 800
rect 396446 0 396502 800
rect 397182 0 397238 800
rect 398010 0 398066 800
rect 398746 0 398802 800
rect 399574 0 399630 800
<< obsm2 >>
rect 1952 399144 4746 399242
rect 4914 399144 7966 399242
rect 8134 399144 11278 399242
rect 11446 399144 14498 399242
rect 14666 399144 17718 399242
rect 17886 399144 21030 399242
rect 21198 399144 24250 399242
rect 24418 399144 27470 399242
rect 27638 399144 30782 399242
rect 30950 399144 34002 399242
rect 34170 399144 37222 399242
rect 37390 399144 40534 399242
rect 40702 399144 43754 399242
rect 43922 399144 46974 399242
rect 47142 399144 50286 399242
rect 50454 399144 53506 399242
rect 53674 399144 56726 399242
rect 56894 399144 60038 399242
rect 60206 399144 63258 399242
rect 63426 399144 66478 399242
rect 66646 399144 69790 399242
rect 69958 399144 73010 399242
rect 73178 399144 76322 399242
rect 76490 399144 79542 399242
rect 79710 399144 82762 399242
rect 82930 399144 86074 399242
rect 86242 399144 89294 399242
rect 89462 399144 92514 399242
rect 92682 399144 95826 399242
rect 95994 399144 99046 399242
rect 99214 399144 102266 399242
rect 102434 399144 105578 399242
rect 105746 399144 108798 399242
rect 108966 399144 112018 399242
rect 112186 399144 115330 399242
rect 115498 399144 118550 399242
rect 118718 399144 121770 399242
rect 121938 399144 125082 399242
rect 125250 399144 128302 399242
rect 128470 399144 131522 399242
rect 131690 399144 134834 399242
rect 135002 399144 138054 399242
rect 138222 399144 141366 399242
rect 141534 399144 144586 399242
rect 144754 399144 147806 399242
rect 147974 399144 151118 399242
rect 151286 399144 154338 399242
rect 154506 399144 157558 399242
rect 157726 399144 160870 399242
rect 161038 399144 164090 399242
rect 164258 399144 167310 399242
rect 167478 399144 170622 399242
rect 170790 399144 173842 399242
rect 174010 399144 177062 399242
rect 177230 399144 180374 399242
rect 180542 399144 183594 399242
rect 183762 399144 186814 399242
rect 186982 399144 190126 399242
rect 190294 399144 193346 399242
rect 193514 399144 196566 399242
rect 196734 399144 199878 399242
rect 200046 399144 203098 399242
rect 203266 399144 206410 399242
rect 206578 399144 209630 399242
rect 209798 399144 212850 399242
rect 213018 399144 216162 399242
rect 216330 399144 219382 399242
rect 219550 399144 222602 399242
rect 222770 399144 225914 399242
rect 226082 399144 229134 399242
rect 229302 399144 232354 399242
rect 232522 399144 235666 399242
rect 235834 399144 238886 399242
rect 239054 399144 242106 399242
rect 242274 399144 245418 399242
rect 245586 399144 248638 399242
rect 248806 399144 251858 399242
rect 252026 399144 255170 399242
rect 255338 399144 258390 399242
rect 258558 399144 261610 399242
rect 261778 399144 264922 399242
rect 265090 399144 268142 399242
rect 268310 399144 271454 399242
rect 271622 399144 274674 399242
rect 274842 399144 277894 399242
rect 278062 399144 281206 399242
rect 281374 399144 284426 399242
rect 284594 399144 287646 399242
rect 287814 399144 290958 399242
rect 291126 399144 294178 399242
rect 294346 399144 297398 399242
rect 297566 399144 300710 399242
rect 300878 399144 303930 399242
rect 304098 399144 307150 399242
rect 307318 399144 310462 399242
rect 310630 399144 313682 399242
rect 313850 399144 316902 399242
rect 317070 399144 320214 399242
rect 320382 399144 323434 399242
rect 323602 399144 326654 399242
rect 326822 399144 329966 399242
rect 330134 399144 333186 399242
rect 333354 399144 336498 399242
rect 336666 399144 339718 399242
rect 339886 399144 342938 399242
rect 343106 399144 346250 399242
rect 346418 399144 349470 399242
rect 349638 399144 352690 399242
rect 352858 399144 356002 399242
rect 356170 399144 359222 399242
rect 359390 399144 362442 399242
rect 362610 399144 365754 399242
rect 365922 399144 368974 399242
rect 369142 399144 372194 399242
rect 372362 399144 375506 399242
rect 375674 399144 378726 399242
rect 378894 399144 381946 399242
rect 382114 399144 385258 399242
rect 385426 399144 388478 399242
rect 388646 399144 389312 399242
rect 1952 856 389312 399144
rect 2062 734 2630 856
rect 2798 734 3458 856
rect 3626 734 4194 856
rect 4362 734 5022 856
rect 5190 734 5850 856
rect 6018 734 6586 856
rect 6754 734 7414 856
rect 7582 734 8150 856
rect 8318 734 8978 856
rect 9146 734 9714 856
rect 9882 734 10542 856
rect 10710 734 11370 856
rect 11538 734 12106 856
rect 12274 734 12934 856
rect 13102 734 13670 856
rect 13838 734 14498 856
rect 14666 734 15234 856
rect 15402 734 16062 856
rect 16230 734 16890 856
rect 17058 734 17626 856
rect 17794 734 18454 856
rect 18622 734 19190 856
rect 19358 734 20018 856
rect 20186 734 20754 856
rect 20922 734 21582 856
rect 21750 734 22410 856
rect 22578 734 23146 856
rect 23314 734 23974 856
rect 24142 734 24710 856
rect 24878 734 25538 856
rect 25706 734 26366 856
rect 26534 734 27102 856
rect 27270 734 27930 856
rect 28098 734 28666 856
rect 28834 734 29494 856
rect 29662 734 30230 856
rect 30398 734 31058 856
rect 31226 734 31886 856
rect 32054 734 32622 856
rect 32790 734 33450 856
rect 33618 734 34186 856
rect 34354 734 35014 856
rect 35182 734 35750 856
rect 35918 734 36578 856
rect 36746 734 37406 856
rect 37574 734 38142 856
rect 38310 734 38970 856
rect 39138 734 39706 856
rect 39874 734 40534 856
rect 40702 734 41270 856
rect 41438 734 42098 856
rect 42266 734 42926 856
rect 43094 734 43662 856
rect 43830 734 44490 856
rect 44658 734 45226 856
rect 45394 734 46054 856
rect 46222 734 46790 856
rect 46958 734 47618 856
rect 47786 734 48446 856
rect 48614 734 49182 856
rect 49350 734 50010 856
rect 50178 734 50746 856
rect 50914 734 51574 856
rect 51742 734 52402 856
rect 52570 734 53138 856
rect 53306 734 53966 856
rect 54134 734 54702 856
rect 54870 734 55530 856
rect 55698 734 56266 856
rect 56434 734 57094 856
rect 57262 734 57922 856
rect 58090 734 58658 856
rect 58826 734 59486 856
rect 59654 734 60222 856
rect 60390 734 61050 856
rect 61218 734 61786 856
rect 61954 734 62614 856
rect 62782 734 63442 856
rect 63610 734 64178 856
rect 64346 734 65006 856
rect 65174 734 65742 856
rect 65910 734 66570 856
rect 66738 734 67306 856
rect 67474 734 68134 856
rect 68302 734 68962 856
rect 69130 734 69698 856
rect 69866 734 70526 856
rect 70694 734 71262 856
rect 71430 734 72090 856
rect 72258 734 72826 856
rect 72994 734 73654 856
rect 73822 734 74482 856
rect 74650 734 75218 856
rect 75386 734 76046 856
rect 76214 734 76782 856
rect 76950 734 77610 856
rect 77778 734 78438 856
rect 78606 734 79174 856
rect 79342 734 80002 856
rect 80170 734 80738 856
rect 80906 734 81566 856
rect 81734 734 82302 856
rect 82470 734 83130 856
rect 83298 734 83958 856
rect 84126 734 84694 856
rect 84862 734 85522 856
rect 85690 734 86258 856
rect 86426 734 87086 856
rect 87254 734 87822 856
rect 87990 734 88650 856
rect 88818 734 89478 856
rect 89646 734 90214 856
rect 90382 734 91042 856
rect 91210 734 91778 856
rect 91946 734 92606 856
rect 92774 734 93342 856
rect 93510 734 94170 856
rect 94338 734 94998 856
rect 95166 734 95734 856
rect 95902 734 96562 856
rect 96730 734 97298 856
rect 97466 734 98126 856
rect 98294 734 98862 856
rect 99030 734 99690 856
rect 99858 734 100518 856
rect 100686 734 101254 856
rect 101422 734 102082 856
rect 102250 734 102818 856
rect 102986 734 103646 856
rect 103814 734 104474 856
rect 104642 734 105210 856
rect 105378 734 106038 856
rect 106206 734 106774 856
rect 106942 734 107602 856
rect 107770 734 108338 856
rect 108506 734 109166 856
rect 109334 734 109994 856
rect 110162 734 110730 856
rect 110898 734 111558 856
rect 111726 734 112294 856
rect 112462 734 113122 856
rect 113290 734 113858 856
rect 114026 734 114686 856
rect 114854 734 115514 856
rect 115682 734 116250 856
rect 116418 734 117078 856
rect 117246 734 117814 856
rect 117982 734 118642 856
rect 118810 734 119378 856
rect 119546 734 120206 856
rect 120374 734 121034 856
rect 121202 734 121770 856
rect 121938 734 122598 856
rect 122766 734 123334 856
rect 123502 734 124162 856
rect 124330 734 124898 856
rect 125066 734 125726 856
rect 125894 734 126554 856
rect 126722 734 127290 856
rect 127458 734 128118 856
rect 128286 734 128854 856
rect 129022 734 129682 856
rect 129850 734 130510 856
rect 130678 734 131246 856
rect 131414 734 132074 856
rect 132242 734 132810 856
rect 132978 734 133638 856
rect 133806 734 134374 856
rect 134542 734 135202 856
rect 135370 734 136030 856
rect 136198 734 136766 856
rect 136934 734 137594 856
rect 137762 734 138330 856
rect 138498 734 139158 856
rect 139326 734 139894 856
rect 140062 734 140722 856
rect 140890 734 141550 856
rect 141718 734 142286 856
rect 142454 734 143114 856
rect 143282 734 143850 856
rect 144018 734 144678 856
rect 144846 734 145414 856
rect 145582 734 146242 856
rect 146410 734 147070 856
rect 147238 734 147806 856
rect 147974 734 148634 856
rect 148802 734 149370 856
rect 149538 734 150198 856
rect 150366 734 151026 856
rect 151194 734 151762 856
rect 151930 734 152590 856
rect 152758 734 153326 856
rect 153494 734 154154 856
rect 154322 734 154890 856
rect 155058 734 155718 856
rect 155886 734 156546 856
rect 156714 734 157282 856
rect 157450 734 158110 856
rect 158278 734 158846 856
rect 159014 734 159674 856
rect 159842 734 160410 856
rect 160578 734 161238 856
rect 161406 734 162066 856
rect 162234 734 162802 856
rect 162970 734 163630 856
rect 163798 734 164366 856
rect 164534 734 165194 856
rect 165362 734 165930 856
rect 166098 734 166758 856
rect 166926 734 167586 856
rect 167754 734 168322 856
rect 168490 734 169150 856
rect 169318 734 169886 856
rect 170054 734 170714 856
rect 170882 734 171450 856
rect 171618 734 172278 856
rect 172446 734 173106 856
rect 173274 734 173842 856
rect 174010 734 174670 856
rect 174838 734 175406 856
rect 175574 734 176234 856
rect 176402 734 177062 856
rect 177230 734 177798 856
rect 177966 734 178626 856
rect 178794 734 179362 856
rect 179530 734 180190 856
rect 180358 734 180926 856
rect 181094 734 181754 856
rect 181922 734 182582 856
rect 182750 734 183318 856
rect 183486 734 184146 856
rect 184314 734 184882 856
rect 185050 734 185710 856
rect 185878 734 186446 856
rect 186614 734 187274 856
rect 187442 734 188102 856
rect 188270 734 188838 856
rect 189006 734 189666 856
rect 189834 734 190402 856
rect 190570 734 191230 856
rect 191398 734 191966 856
rect 192134 734 192794 856
rect 192962 734 193622 856
rect 193790 734 194358 856
rect 194526 734 195186 856
rect 195354 734 195922 856
rect 196090 734 196750 856
rect 196918 734 197486 856
rect 197654 734 198314 856
rect 198482 734 199142 856
rect 199310 734 199878 856
rect 200046 734 200706 856
rect 200874 734 201442 856
rect 201610 734 202270 856
rect 202438 734 203098 856
rect 203266 734 203834 856
rect 204002 734 204662 856
rect 204830 734 205398 856
rect 205566 734 206226 856
rect 206394 734 206962 856
rect 207130 734 207790 856
rect 207958 734 208618 856
rect 208786 734 209354 856
rect 209522 734 210182 856
rect 210350 734 210918 856
rect 211086 734 211746 856
rect 211914 734 212482 856
rect 212650 734 213310 856
rect 213478 734 214138 856
rect 214306 734 214874 856
rect 215042 734 215702 856
rect 215870 734 216438 856
rect 216606 734 217266 856
rect 217434 734 218002 856
rect 218170 734 218830 856
rect 218998 734 219658 856
rect 219826 734 220394 856
rect 220562 734 221222 856
rect 221390 734 221958 856
rect 222126 734 222786 856
rect 222954 734 223522 856
rect 223690 734 224350 856
rect 224518 734 225178 856
rect 225346 734 225914 856
rect 226082 734 226742 856
rect 226910 734 227478 856
rect 227646 734 228306 856
rect 228474 734 229134 856
rect 229302 734 229870 856
rect 230038 734 230698 856
rect 230866 734 231434 856
rect 231602 734 232262 856
rect 232430 734 232998 856
rect 233166 734 233826 856
rect 233994 734 234654 856
rect 234822 734 235390 856
rect 235558 734 236218 856
rect 236386 734 236954 856
rect 237122 734 237782 856
rect 237950 734 238518 856
rect 238686 734 239346 856
rect 239514 734 240174 856
rect 240342 734 240910 856
rect 241078 734 241738 856
rect 241906 734 242474 856
rect 242642 734 243302 856
rect 243470 734 244038 856
rect 244206 734 244866 856
rect 245034 734 245694 856
rect 245862 734 246430 856
rect 246598 734 247258 856
rect 247426 734 247994 856
rect 248162 734 248822 856
rect 248990 734 249558 856
rect 249726 734 250386 856
rect 250554 734 251214 856
rect 251382 734 251950 856
rect 252118 734 252778 856
rect 252946 734 253514 856
rect 253682 734 254342 856
rect 254510 734 255170 856
rect 255338 734 255906 856
rect 256074 734 256734 856
rect 256902 734 257470 856
rect 257638 734 258298 856
rect 258466 734 259034 856
rect 259202 734 259862 856
rect 260030 734 260690 856
rect 260858 734 261426 856
rect 261594 734 262254 856
rect 262422 734 262990 856
rect 263158 734 263818 856
rect 263986 734 264554 856
rect 264722 734 265382 856
rect 265550 734 266210 856
rect 266378 734 266946 856
rect 267114 734 267774 856
rect 267942 734 268510 856
rect 268678 734 269338 856
rect 269506 734 270074 856
rect 270242 734 270902 856
rect 271070 734 271730 856
rect 271898 734 272466 856
rect 272634 734 273294 856
rect 273462 734 274030 856
rect 274198 734 274858 856
rect 275026 734 275686 856
rect 275854 734 276422 856
rect 276590 734 277250 856
rect 277418 734 277986 856
rect 278154 734 278814 856
rect 278982 734 279550 856
rect 279718 734 280378 856
rect 280546 734 281206 856
rect 281374 734 281942 856
rect 282110 734 282770 856
rect 282938 734 283506 856
rect 283674 734 284334 856
rect 284502 734 285070 856
rect 285238 734 285898 856
rect 286066 734 286726 856
rect 286894 734 287462 856
rect 287630 734 288290 856
rect 288458 734 289026 856
rect 289194 734 289854 856
rect 290022 734 290590 856
rect 290758 734 291418 856
rect 291586 734 292246 856
rect 292414 734 292982 856
rect 293150 734 293810 856
rect 293978 734 294546 856
rect 294714 734 295374 856
rect 295542 734 296110 856
rect 296278 734 296938 856
rect 297106 734 297766 856
rect 297934 734 298502 856
rect 298670 734 299330 856
rect 299498 734 300066 856
rect 300234 734 300894 856
rect 301062 734 301722 856
rect 301890 734 302458 856
rect 302626 734 303286 856
rect 303454 734 304022 856
rect 304190 734 304850 856
rect 305018 734 305586 856
rect 305754 734 306414 856
rect 306582 734 307242 856
rect 307410 734 307978 856
rect 308146 734 308806 856
rect 308974 734 309542 856
rect 309710 734 310370 856
rect 310538 734 311106 856
rect 311274 734 311934 856
rect 312102 734 312762 856
rect 312930 734 313498 856
rect 313666 734 314326 856
rect 314494 734 315062 856
rect 315230 734 315890 856
rect 316058 734 316626 856
rect 316794 734 317454 856
rect 317622 734 318282 856
rect 318450 734 319018 856
rect 319186 734 319846 856
rect 320014 734 320582 856
rect 320750 734 321410 856
rect 321578 734 322146 856
rect 322314 734 322974 856
rect 323142 734 323802 856
rect 323970 734 324538 856
rect 324706 734 325366 856
rect 325534 734 326102 856
rect 326270 734 326930 856
rect 327098 734 327758 856
rect 327926 734 328494 856
rect 328662 734 329322 856
rect 329490 734 330058 856
rect 330226 734 330886 856
rect 331054 734 331622 856
rect 331790 734 332450 856
rect 332618 734 333278 856
rect 333446 734 334014 856
rect 334182 734 334842 856
rect 335010 734 335578 856
rect 335746 734 336406 856
rect 336574 734 337142 856
rect 337310 734 337970 856
rect 338138 734 338798 856
rect 338966 734 339534 856
rect 339702 734 340362 856
rect 340530 734 341098 856
rect 341266 734 341926 856
rect 342094 734 342662 856
rect 342830 734 343490 856
rect 343658 734 344318 856
rect 344486 734 345054 856
rect 345222 734 345882 856
rect 346050 734 346618 856
rect 346786 734 347446 856
rect 347614 734 348182 856
rect 348350 734 349010 856
rect 349178 734 349838 856
rect 350006 734 350574 856
rect 350742 734 351402 856
rect 351570 734 352138 856
rect 352306 734 352966 856
rect 353134 734 353794 856
rect 353962 734 354530 856
rect 354698 734 355358 856
rect 355526 734 356094 856
rect 356262 734 356922 856
rect 357090 734 357658 856
rect 357826 734 358486 856
rect 358654 734 359314 856
rect 359482 734 360050 856
rect 360218 734 360878 856
rect 361046 734 361614 856
rect 361782 734 362442 856
rect 362610 734 363178 856
rect 363346 734 364006 856
rect 364174 734 364834 856
rect 365002 734 365570 856
rect 365738 734 366398 856
rect 366566 734 367134 856
rect 367302 734 367962 856
rect 368130 734 368698 856
rect 368866 734 369526 856
rect 369694 734 370354 856
rect 370522 734 371090 856
rect 371258 734 371918 856
rect 372086 734 372654 856
rect 372822 734 373482 856
rect 373650 734 374218 856
rect 374386 734 375046 856
rect 375214 734 375874 856
rect 376042 734 376610 856
rect 376778 734 377438 856
rect 377606 734 378174 856
rect 378342 734 379002 856
rect 379170 734 379830 856
rect 379998 734 380566 856
rect 380734 734 381394 856
rect 381562 734 382130 856
rect 382298 734 382958 856
rect 383126 734 383694 856
rect 383862 734 384522 856
rect 384690 734 385350 856
rect 385518 734 386086 856
rect 386254 734 386914 856
rect 387082 734 387650 856
rect 387818 734 388478 856
rect 388646 734 389214 856
<< metal3 >>
rect 0 333208 800 333328
rect 0 199928 800 200048
rect 0 66648 800 66768
rect 399200 349800 400000 349920
rect 399200 249840 400000 249960
rect 399200 149880 400000 150000
rect 399200 49920 400000 50040
<< obsm3 >>
rect 4208 2143 388528 397697
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
rect 203888 2128 204208 397712
rect 219248 2128 219568 397712
rect 234608 2128 234928 397712
rect 249968 2128 250288 397712
rect 265328 2128 265648 397712
rect 280688 2128 281008 397712
rect 296048 2128 296368 397712
rect 311408 2128 311728 397712
rect 326768 2128 327088 397712
rect 342128 2128 342448 397712
rect 357488 2128 357808 397712
rect 372848 2128 373168 397712
rect 388208 2128 388528 397712
<< obsm4 >>
rect 55443 21659 65568 397357
rect 66048 21659 80928 397357
rect 81408 21659 96288 397357
rect 96768 21659 111648 397357
rect 112128 21659 127008 397357
rect 127488 21659 142368 397357
rect 142848 21659 157728 397357
rect 158208 21659 173088 397357
rect 173568 21659 188448 397357
rect 188928 21659 203808 397357
rect 204288 21659 219168 397357
rect 219648 21659 234528 397357
rect 235008 21659 249888 397357
rect 250368 21659 265248 397357
rect 265728 21659 280608 397357
rect 281088 21659 295813 397357
<< labels >>
rlabel metal2 s 390098 0 390154 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 66648 800 66768 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 385314 399200 385370 400000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 394054 0 394110 800 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 394790 0 394846 800 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 399200 149880 400000 150000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 395618 0 395674 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 396446 0 396502 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 388534 399200 388590 400000 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 397182 0 397238 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 199928 800 200048 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 390926 0 390982 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 391754 399200 391810 400000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 398010 0 398066 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 395066 399200 395122 400000 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 399200 249840 400000 249960 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 398286 399200 398342 400000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 398746 0 398802 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 333208 800 333328 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 399200 349800 400000 349920 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 399574 0 399630 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 391662 0 391718 800 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal2 s 372250 399200 372306 400000 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 392490 0 392546 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal2 s 375562 399200 375618 400000 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 399200 49920 400000 50040 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 378782 399200 378838 400000 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 382002 399200 382058 400000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 393226 0 393282 800 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 1582 399200 1638 400000 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 99102 399200 99158 400000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 108854 399200 108910 400000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 118606 399200 118662 400000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 128358 399200 128414 400000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 138110 399200 138166 400000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 147862 399200 147918 400000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 157614 399200 157670 400000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 167366 399200 167422 400000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 177118 399200 177174 400000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 186870 399200 186926 400000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 11334 399200 11390 400000 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 196622 399200 196678 400000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 206466 399200 206522 400000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 216218 399200 216274 400000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 225970 399200 226026 400000 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 235722 399200 235778 400000 6 io_in[24]
port 46 nsew signal input
rlabel metal2 s 245474 399200 245530 400000 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 255226 399200 255282 400000 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 264978 399200 265034 400000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 274730 399200 274786 400000 6 io_in[28]
port 50 nsew signal input
rlabel metal2 s 284482 399200 284538 400000 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 21086 399200 21142 400000 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 294234 399200 294290 400000 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 303986 399200 304042 400000 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 313738 399200 313794 400000 6 io_in[32]
port 55 nsew signal input
rlabel metal2 s 323490 399200 323546 400000 6 io_in[33]
port 56 nsew signal input
rlabel metal2 s 333242 399200 333298 400000 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 342994 399200 343050 400000 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 352746 399200 352802 400000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 362498 399200 362554 400000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 30838 399200 30894 400000 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 40590 399200 40646 400000 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 50342 399200 50398 400000 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 60094 399200 60150 400000 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 69846 399200 69902 400000 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 79598 399200 79654 400000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 89350 399200 89406 400000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 4802 399200 4858 400000 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 102322 399200 102378 400000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 112074 399200 112130 400000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 121826 399200 121882 400000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 131578 399200 131634 400000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 141422 399200 141478 400000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 151174 399200 151230 400000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 160926 399200 160982 400000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 170678 399200 170734 400000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 180430 399200 180486 400000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 190182 399200 190238 400000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 14554 399200 14610 400000 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 199934 399200 199990 400000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 209686 399200 209742 400000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 219438 399200 219494 400000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 229190 399200 229246 400000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal2 s 238942 399200 238998 400000 6 io_oeb[24]
port 84 nsew signal output
rlabel metal2 s 248694 399200 248750 400000 6 io_oeb[25]
port 85 nsew signal output
rlabel metal2 s 258446 399200 258502 400000 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 268198 399200 268254 400000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 277950 399200 278006 400000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal2 s 287702 399200 287758 400000 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 24306 399200 24362 400000 6 io_oeb[2]
port 90 nsew signal output
rlabel metal2 s 297454 399200 297510 400000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 307206 399200 307262 400000 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 316958 399200 317014 400000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal2 s 326710 399200 326766 400000 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 336554 399200 336610 400000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 346306 399200 346362 400000 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 356058 399200 356114 400000 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 365810 399200 365866 400000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 34058 399200 34114 400000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 43810 399200 43866 400000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 53562 399200 53618 400000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 63314 399200 63370 400000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 73066 399200 73122 400000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 82818 399200 82874 400000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 92570 399200 92626 400000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 8022 399200 8078 400000 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 105634 399200 105690 400000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 115386 399200 115442 400000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 125138 399200 125194 400000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 134890 399200 134946 400000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 144642 399200 144698 400000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 154394 399200 154450 400000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 164146 399200 164202 400000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 173898 399200 173954 400000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 183650 399200 183706 400000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 193402 399200 193458 400000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 17774 399200 17830 400000 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 203154 399200 203210 400000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 212906 399200 212962 400000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 222658 399200 222714 400000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 232410 399200 232466 400000 6 io_out[23]
port 121 nsew signal output
rlabel metal2 s 242162 399200 242218 400000 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 251914 399200 251970 400000 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 261666 399200 261722 400000 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 271510 399200 271566 400000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 281262 399200 281318 400000 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 291014 399200 291070 400000 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 27526 399200 27582 400000 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 300766 399200 300822 400000 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 310518 399200 310574 400000 6 io_out[31]
port 130 nsew signal output
rlabel metal2 s 320270 399200 320326 400000 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 330022 399200 330078 400000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 339774 399200 339830 400000 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 349526 399200 349582 400000 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 359278 399200 359334 400000 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 369030 399200 369086 400000 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 37278 399200 37334 400000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 47030 399200 47086 400000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 56782 399200 56838 400000 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 66534 399200 66590 400000 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 76378 399200 76434 400000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 86130 399200 86186 400000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 95882 399200 95938 400000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 386970 0 387026 800 6 irq[0]
port 144 nsew signal output
rlabel metal2 s 387706 0 387762 800 6 irq[1]
port 145 nsew signal output
rlabel metal2 s 388534 0 388590 800 6 irq[2]
port 146 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 la_data_in[0]
port 147 nsew signal input
rlabel metal2 s 320638 0 320694 800 6 la_data_in[100]
port 148 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 la_data_in[101]
port 149 nsew signal input
rlabel metal2 s 325422 0 325478 800 6 la_data_in[102]
port 150 nsew signal input
rlabel metal2 s 327814 0 327870 800 6 la_data_in[103]
port 151 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[104]
port 152 nsew signal input
rlabel metal2 s 332506 0 332562 800 6 la_data_in[105]
port 153 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 la_data_in[106]
port 154 nsew signal input
rlabel metal2 s 337198 0 337254 800 6 la_data_in[107]
port 155 nsew signal input
rlabel metal2 s 339590 0 339646 800 6 la_data_in[108]
port 156 nsew signal input
rlabel metal2 s 341982 0 342038 800 6 la_data_in[109]
port 157 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[10]
port 158 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_data_in[110]
port 159 nsew signal input
rlabel metal2 s 346674 0 346730 800 6 la_data_in[111]
port 160 nsew signal input
rlabel metal2 s 349066 0 349122 800 6 la_data_in[112]
port 161 nsew signal input
rlabel metal2 s 351458 0 351514 800 6 la_data_in[113]
port 162 nsew signal input
rlabel metal2 s 353850 0 353906 800 6 la_data_in[114]
port 163 nsew signal input
rlabel metal2 s 356150 0 356206 800 6 la_data_in[115]
port 164 nsew signal input
rlabel metal2 s 358542 0 358598 800 6 la_data_in[116]
port 165 nsew signal input
rlabel metal2 s 360934 0 360990 800 6 la_data_in[117]
port 166 nsew signal input
rlabel metal2 s 363234 0 363290 800 6 la_data_in[118]
port 167 nsew signal input
rlabel metal2 s 365626 0 365682 800 6 la_data_in[119]
port 168 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_data_in[11]
port 169 nsew signal input
rlabel metal2 s 368018 0 368074 800 6 la_data_in[120]
port 170 nsew signal input
rlabel metal2 s 370410 0 370466 800 6 la_data_in[121]
port 171 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_data_in[122]
port 172 nsew signal input
rlabel metal2 s 375102 0 375158 800 6 la_data_in[123]
port 173 nsew signal input
rlabel metal2 s 377494 0 377550 800 6 la_data_in[124]
port 174 nsew signal input
rlabel metal2 s 379886 0 379942 800 6 la_data_in[125]
port 175 nsew signal input
rlabel metal2 s 382186 0 382242 800 6 la_data_in[126]
port 176 nsew signal input
rlabel metal2 s 384578 0 384634 800 6 la_data_in[127]
port 177 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[12]
port 178 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[13]
port 179 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[14]
port 180 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[15]
port 181 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[16]
port 182 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[17]
port 183 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_data_in[18]
port 184 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[19]
port 185 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[1]
port 186 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[20]
port 187 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_data_in[21]
port 188 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_data_in[22]
port 189 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[23]
port 190 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[24]
port 191 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[25]
port 192 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[26]
port 193 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[27]
port 194 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[28]
port 195 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_data_in[29]
port 196 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[2]
port 197 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[30]
port 198 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[31]
port 199 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[32]
port 200 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[33]
port 201 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[34]
port 202 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[35]
port 203 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_data_in[36]
port 204 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[37]
port 205 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_data_in[38]
port 206 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_data_in[39]
port 207 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[3]
port 208 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[40]
port 209 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[41]
port 210 nsew signal input
rlabel metal2 s 183374 0 183430 800 6 la_data_in[42]
port 211 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_data_in[43]
port 212 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[44]
port 213 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_data_in[45]
port 214 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_data_in[46]
port 215 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[47]
port 216 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[48]
port 217 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[49]
port 218 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[4]
port 219 nsew signal input
rlabel metal2 s 202326 0 202382 800 6 la_data_in[50]
port 220 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[51]
port 221 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_data_in[52]
port 222 nsew signal input
rlabel metal2 s 209410 0 209466 800 6 la_data_in[53]
port 223 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[54]
port 224 nsew signal input
rlabel metal2 s 214194 0 214250 800 6 la_data_in[55]
port 225 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[56]
port 226 nsew signal input
rlabel metal2 s 218886 0 218942 800 6 la_data_in[57]
port 227 nsew signal input
rlabel metal2 s 221278 0 221334 800 6 la_data_in[58]
port 228 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_data_in[59]
port 229 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[5]
port 230 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_data_in[60]
port 231 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[61]
port 232 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_data_in[62]
port 233 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_data_in[63]
port 234 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_data_in[64]
port 235 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[65]
port 236 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[66]
port 237 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_data_in[67]
port 238 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_data_in[68]
port 239 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_data_in[69]
port 240 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[6]
port 241 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_data_in[70]
port 242 nsew signal input
rlabel metal2 s 252006 0 252062 800 6 la_data_in[71]
port 243 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[72]
port 244 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_data_in[73]
port 245 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 la_data_in[74]
port 246 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 la_data_in[75]
port 247 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_data_in[76]
port 248 nsew signal input
rlabel metal2 s 266266 0 266322 800 6 la_data_in[77]
port 249 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 la_data_in[78]
port 250 nsew signal input
rlabel metal2 s 270958 0 271014 800 6 la_data_in[79]
port 251 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[7]
port 252 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_data_in[80]
port 253 nsew signal input
rlabel metal2 s 275742 0 275798 800 6 la_data_in[81]
port 254 nsew signal input
rlabel metal2 s 278042 0 278098 800 6 la_data_in[82]
port 255 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_data_in[83]
port 256 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[84]
port 257 nsew signal input
rlabel metal2 s 285126 0 285182 800 6 la_data_in[85]
port 258 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_data_in[86]
port 259 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 la_data_in[87]
port 260 nsew signal input
rlabel metal2 s 292302 0 292358 800 6 la_data_in[88]
port 261 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_data_in[89]
port 262 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_data_in[8]
port 263 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_data_in[90]
port 264 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_data_in[91]
port 265 nsew signal input
rlabel metal2 s 301778 0 301834 800 6 la_data_in[92]
port 266 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_data_in[93]
port 267 nsew signal input
rlabel metal2 s 306470 0 306526 800 6 la_data_in[94]
port 268 nsew signal input
rlabel metal2 s 308862 0 308918 800 6 la_data_in[95]
port 269 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 la_data_in[96]
port 270 nsew signal input
rlabel metal2 s 313554 0 313610 800 6 la_data_in[97]
port 271 nsew signal input
rlabel metal2 s 315946 0 316002 800 6 la_data_in[98]
port 272 nsew signal input
rlabel metal2 s 318338 0 318394 800 6 la_data_in[99]
port 273 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[9]
port 274 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_out[0]
port 275 nsew signal output
rlabel metal2 s 321466 0 321522 800 6 la_data_out[100]
port 276 nsew signal output
rlabel metal2 s 323858 0 323914 800 6 la_data_out[101]
port 277 nsew signal output
rlabel metal2 s 326158 0 326214 800 6 la_data_out[102]
port 278 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 la_data_out[103]
port 279 nsew signal output
rlabel metal2 s 330942 0 330998 800 6 la_data_out[104]
port 280 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[105]
port 281 nsew signal output
rlabel metal2 s 335634 0 335690 800 6 la_data_out[106]
port 282 nsew signal output
rlabel metal2 s 338026 0 338082 800 6 la_data_out[107]
port 283 nsew signal output
rlabel metal2 s 340418 0 340474 800 6 la_data_out[108]
port 284 nsew signal output
rlabel metal2 s 342718 0 342774 800 6 la_data_out[109]
port 285 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[10]
port 286 nsew signal output
rlabel metal2 s 345110 0 345166 800 6 la_data_out[110]
port 287 nsew signal output
rlabel metal2 s 347502 0 347558 800 6 la_data_out[111]
port 288 nsew signal output
rlabel metal2 s 349894 0 349950 800 6 la_data_out[112]
port 289 nsew signal output
rlabel metal2 s 352194 0 352250 800 6 la_data_out[113]
port 290 nsew signal output
rlabel metal2 s 354586 0 354642 800 6 la_data_out[114]
port 291 nsew signal output
rlabel metal2 s 356978 0 357034 800 6 la_data_out[115]
port 292 nsew signal output
rlabel metal2 s 359370 0 359426 800 6 la_data_out[116]
port 293 nsew signal output
rlabel metal2 s 361670 0 361726 800 6 la_data_out[117]
port 294 nsew signal output
rlabel metal2 s 364062 0 364118 800 6 la_data_out[118]
port 295 nsew signal output
rlabel metal2 s 366454 0 366510 800 6 la_data_out[119]
port 296 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[11]
port 297 nsew signal output
rlabel metal2 s 368754 0 368810 800 6 la_data_out[120]
port 298 nsew signal output
rlabel metal2 s 371146 0 371202 800 6 la_data_out[121]
port 299 nsew signal output
rlabel metal2 s 373538 0 373594 800 6 la_data_out[122]
port 300 nsew signal output
rlabel metal2 s 375930 0 375986 800 6 la_data_out[123]
port 301 nsew signal output
rlabel metal2 s 378230 0 378286 800 6 la_data_out[124]
port 302 nsew signal output
rlabel metal2 s 380622 0 380678 800 6 la_data_out[125]
port 303 nsew signal output
rlabel metal2 s 383014 0 383070 800 6 la_data_out[126]
port 304 nsew signal output
rlabel metal2 s 385406 0 385462 800 6 la_data_out[127]
port 305 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[12]
port 306 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[13]
port 307 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[14]
port 308 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 la_data_out[15]
port 309 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[16]
port 310 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[17]
port 311 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[18]
port 312 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[19]
port 313 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[1]
port 314 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[20]
port 315 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[21]
port 316 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[22]
port 317 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[23]
port 318 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[24]
port 319 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[25]
port 320 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[26]
port 321 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[27]
port 322 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[28]
port 323 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[29]
port 324 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[2]
port 325 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[30]
port 326 nsew signal output
rlabel metal2 s 158166 0 158222 800 6 la_data_out[31]
port 327 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[32]
port 328 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[33]
port 329 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 la_data_out[34]
port 330 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[35]
port 331 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[36]
port 332 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[37]
port 333 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[38]
port 334 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 la_data_out[39]
port 335 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[3]
port 336 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[40]
port 337 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[41]
port 338 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[42]
port 339 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[43]
port 340 nsew signal output
rlabel metal2 s 188894 0 188950 800 6 la_data_out[44]
port 341 nsew signal output
rlabel metal2 s 191286 0 191342 800 6 la_data_out[45]
port 342 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 la_data_out[46]
port 343 nsew signal output
rlabel metal2 s 195978 0 196034 800 6 la_data_out[47]
port 344 nsew signal output
rlabel metal2 s 198370 0 198426 800 6 la_data_out[48]
port 345 nsew signal output
rlabel metal2 s 200762 0 200818 800 6 la_data_out[49]
port 346 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[4]
port 347 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 la_data_out[50]
port 348 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[51]
port 349 nsew signal output
rlabel metal2 s 207846 0 207902 800 6 la_data_out[52]
port 350 nsew signal output
rlabel metal2 s 210238 0 210294 800 6 la_data_out[53]
port 351 nsew signal output
rlabel metal2 s 212538 0 212594 800 6 la_data_out[54]
port 352 nsew signal output
rlabel metal2 s 214930 0 214986 800 6 la_data_out[55]
port 353 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 la_data_out[56]
port 354 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 la_data_out[57]
port 355 nsew signal output
rlabel metal2 s 222014 0 222070 800 6 la_data_out[58]
port 356 nsew signal output
rlabel metal2 s 224406 0 224462 800 6 la_data_out[59]
port 357 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[5]
port 358 nsew signal output
rlabel metal2 s 226798 0 226854 800 6 la_data_out[60]
port 359 nsew signal output
rlabel metal2 s 229190 0 229246 800 6 la_data_out[61]
port 360 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[62]
port 361 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[63]
port 362 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[64]
port 363 nsew signal output
rlabel metal2 s 238574 0 238630 800 6 la_data_out[65]
port 364 nsew signal output
rlabel metal2 s 240966 0 241022 800 6 la_data_out[66]
port 365 nsew signal output
rlabel metal2 s 243358 0 243414 800 6 la_data_out[67]
port 366 nsew signal output
rlabel metal2 s 245750 0 245806 800 6 la_data_out[68]
port 367 nsew signal output
rlabel metal2 s 248050 0 248106 800 6 la_data_out[69]
port 368 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[6]
port 369 nsew signal output
rlabel metal2 s 250442 0 250498 800 6 la_data_out[70]
port 370 nsew signal output
rlabel metal2 s 252834 0 252890 800 6 la_data_out[71]
port 371 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[72]
port 372 nsew signal output
rlabel metal2 s 257526 0 257582 800 6 la_data_out[73]
port 373 nsew signal output
rlabel metal2 s 259918 0 259974 800 6 la_data_out[74]
port 374 nsew signal output
rlabel metal2 s 262310 0 262366 800 6 la_data_out[75]
port 375 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[76]
port 376 nsew signal output
rlabel metal2 s 267002 0 267058 800 6 la_data_out[77]
port 377 nsew signal output
rlabel metal2 s 269394 0 269450 800 6 la_data_out[78]
port 378 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 la_data_out[79]
port 379 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[7]
port 380 nsew signal output
rlabel metal2 s 274086 0 274142 800 6 la_data_out[80]
port 381 nsew signal output
rlabel metal2 s 276478 0 276534 800 6 la_data_out[81]
port 382 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 la_data_out[82]
port 383 nsew signal output
rlabel metal2 s 281262 0 281318 800 6 la_data_out[83]
port 384 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 la_data_out[84]
port 385 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[85]
port 386 nsew signal output
rlabel metal2 s 288346 0 288402 800 6 la_data_out[86]
port 387 nsew signal output
rlabel metal2 s 290646 0 290702 800 6 la_data_out[87]
port 388 nsew signal output
rlabel metal2 s 293038 0 293094 800 6 la_data_out[88]
port 389 nsew signal output
rlabel metal2 s 295430 0 295486 800 6 la_data_out[89]
port 390 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[8]
port 391 nsew signal output
rlabel metal2 s 297822 0 297878 800 6 la_data_out[90]
port 392 nsew signal output
rlabel metal2 s 300122 0 300178 800 6 la_data_out[91]
port 393 nsew signal output
rlabel metal2 s 302514 0 302570 800 6 la_data_out[92]
port 394 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[93]
port 395 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 la_data_out[94]
port 396 nsew signal output
rlabel metal2 s 309598 0 309654 800 6 la_data_out[95]
port 397 nsew signal output
rlabel metal2 s 311990 0 312046 800 6 la_data_out[96]
port 398 nsew signal output
rlabel metal2 s 314382 0 314438 800 6 la_data_out[97]
port 399 nsew signal output
rlabel metal2 s 316682 0 316738 800 6 la_data_out[98]
port 400 nsew signal output
rlabel metal2 s 319074 0 319130 800 6 la_data_out[99]
port 401 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 la_data_out[9]
port 402 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_oenb[0]
port 403 nsew signal input
rlabel metal2 s 322202 0 322258 800 6 la_oenb[100]
port 404 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 la_oenb[101]
port 405 nsew signal input
rlabel metal2 s 326986 0 327042 800 6 la_oenb[102]
port 406 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_oenb[103]
port 407 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_oenb[104]
port 408 nsew signal input
rlabel metal2 s 334070 0 334126 800 6 la_oenb[105]
port 409 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[106]
port 410 nsew signal input
rlabel metal2 s 338854 0 338910 800 6 la_oenb[107]
port 411 nsew signal input
rlabel metal2 s 341154 0 341210 800 6 la_oenb[108]
port 412 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_oenb[109]
port 413 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[10]
port 414 nsew signal input
rlabel metal2 s 345938 0 345994 800 6 la_oenb[110]
port 415 nsew signal input
rlabel metal2 s 348238 0 348294 800 6 la_oenb[111]
port 416 nsew signal input
rlabel metal2 s 350630 0 350686 800 6 la_oenb[112]
port 417 nsew signal input
rlabel metal2 s 353022 0 353078 800 6 la_oenb[113]
port 418 nsew signal input
rlabel metal2 s 355414 0 355470 800 6 la_oenb[114]
port 419 nsew signal input
rlabel metal2 s 357714 0 357770 800 6 la_oenb[115]
port 420 nsew signal input
rlabel metal2 s 360106 0 360162 800 6 la_oenb[116]
port 421 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 la_oenb[117]
port 422 nsew signal input
rlabel metal2 s 364890 0 364946 800 6 la_oenb[118]
port 423 nsew signal input
rlabel metal2 s 367190 0 367246 800 6 la_oenb[119]
port 424 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[11]
port 425 nsew signal input
rlabel metal2 s 369582 0 369638 800 6 la_oenb[120]
port 426 nsew signal input
rlabel metal2 s 371974 0 372030 800 6 la_oenb[121]
port 427 nsew signal input
rlabel metal2 s 374274 0 374330 800 6 la_oenb[122]
port 428 nsew signal input
rlabel metal2 s 376666 0 376722 800 6 la_oenb[123]
port 429 nsew signal input
rlabel metal2 s 379058 0 379114 800 6 la_oenb[124]
port 430 nsew signal input
rlabel metal2 s 381450 0 381506 800 6 la_oenb[125]
port 431 nsew signal input
rlabel metal2 s 383750 0 383806 800 6 la_oenb[126]
port 432 nsew signal input
rlabel metal2 s 386142 0 386198 800 6 la_oenb[127]
port 433 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[12]
port 434 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[13]
port 435 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[14]
port 436 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[15]
port 437 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[16]
port 438 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[17]
port 439 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[18]
port 440 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[19]
port 441 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[1]
port 442 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_oenb[20]
port 443 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[21]
port 444 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_oenb[22]
port 445 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[23]
port 446 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[24]
port 447 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[25]
port 448 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[26]
port 449 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[27]
port 450 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_oenb[28]
port 451 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[29]
port 452 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[2]
port 453 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[30]
port 454 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[31]
port 455 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_oenb[32]
port 456 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[33]
port 457 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_oenb[34]
port 458 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[35]
port 459 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[36]
port 460 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oenb[37]
port 461 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[38]
port 462 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oenb[39]
port 463 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[3]
port 464 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[40]
port 465 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[41]
port 466 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[42]
port 467 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 la_oenb[43]
port 468 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_oenb[44]
port 469 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[45]
port 470 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oenb[46]
port 471 nsew signal input
rlabel metal2 s 196806 0 196862 800 6 la_oenb[47]
port 472 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[48]
port 473 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_oenb[49]
port 474 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[4]
port 475 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 la_oenb[50]
port 476 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_oenb[51]
port 477 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_oenb[52]
port 478 nsew signal input
rlabel metal2 s 210974 0 211030 800 6 la_oenb[53]
port 479 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_oenb[54]
port 480 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_oenb[55]
port 481 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[56]
port 482 nsew signal input
rlabel metal2 s 220450 0 220506 800 6 la_oenb[57]
port 483 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_oenb[58]
port 484 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oenb[59]
port 485 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_oenb[5]
port 486 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_oenb[60]
port 487 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[61]
port 488 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[62]
port 489 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_oenb[63]
port 490 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_oenb[64]
port 491 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_oenb[65]
port 492 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[66]
port 493 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_oenb[67]
port 494 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_oenb[68]
port 495 nsew signal input
rlabel metal2 s 248878 0 248934 800 6 la_oenb[69]
port 496 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[6]
port 497 nsew signal input
rlabel metal2 s 251270 0 251326 800 6 la_oenb[70]
port 498 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_oenb[71]
port 499 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_oenb[72]
port 500 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oenb[73]
port 501 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_oenb[74]
port 502 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[75]
port 503 nsew signal input
rlabel metal2 s 265438 0 265494 800 6 la_oenb[76]
port 504 nsew signal input
rlabel metal2 s 267830 0 267886 800 6 la_oenb[77]
port 505 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_oenb[78]
port 506 nsew signal input
rlabel metal2 s 272522 0 272578 800 6 la_oenb[79]
port 507 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_oenb[7]
port 508 nsew signal input
rlabel metal2 s 274914 0 274970 800 6 la_oenb[80]
port 509 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 la_oenb[81]
port 510 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_oenb[82]
port 511 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[83]
port 512 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 la_oenb[84]
port 513 nsew signal input
rlabel metal2 s 286782 0 286838 800 6 la_oenb[85]
port 514 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_oenb[86]
port 515 nsew signal input
rlabel metal2 s 291474 0 291530 800 6 la_oenb[87]
port 516 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_oenb[88]
port 517 nsew signal input
rlabel metal2 s 296166 0 296222 800 6 la_oenb[89]
port 518 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_oenb[8]
port 519 nsew signal input
rlabel metal2 s 298558 0 298614 800 6 la_oenb[90]
port 520 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_oenb[91]
port 521 nsew signal input
rlabel metal2 s 303342 0 303398 800 6 la_oenb[92]
port 522 nsew signal input
rlabel metal2 s 305642 0 305698 800 6 la_oenb[93]
port 523 nsew signal input
rlabel metal2 s 308034 0 308090 800 6 la_oenb[94]
port 524 nsew signal input
rlabel metal2 s 310426 0 310482 800 6 la_oenb[95]
port 525 nsew signal input
rlabel metal2 s 312818 0 312874 800 6 la_oenb[96]
port 526 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_oenb[97]
port 527 nsew signal input
rlabel metal2 s 317510 0 317566 800 6 la_oenb[98]
port 528 nsew signal input
rlabel metal2 s 319902 0 319958 800 6 la_oenb[99]
port 529 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[9]
port 530 nsew signal input
rlabel metal2 s 389270 0 389326 800 6 user_clock2
port 531 nsew signal input
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 219248 2128 219568 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 249968 2128 250288 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 280688 2128 281008 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 311408 2128 311728 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 342128 2128 342448 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 372848 2128 373168 397712 6 vccd1
port 532 nsew power input
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 203888 2128 204208 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 234608 2128 234928 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 265328 2128 265648 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 296048 2128 296368 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 326768 2128 327088 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 357488 2128 357808 397712 6 vssd1
port 533 nsew ground input
rlabel metal4 s 388208 2128 388528 397712 6 vssd1
port 533 nsew ground input
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 400000
string LEFview TRUE
string GDS_FILE /home/harald/caravel_mpw5/iic-audiodac-v1/openlane/user_proj_dac/runs/user_proj_dac/results/magic/user_proj_dac.gds
string GDS_END 196621218
string GDS_START 987988
<< end >>

