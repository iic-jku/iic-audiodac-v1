magic
tech sky130A
magscale 1 2
timestamp 1644674034
<< nwell >>
rect 1066 397381 198850 397702
rect 1066 396293 198850 396859
rect 1066 395205 198850 395771
rect 1066 394117 198850 394683
rect 1066 393029 198850 393595
rect 1066 391941 198850 392507
rect 1066 390853 198850 391419
rect 1066 389765 198850 390331
rect 1066 388677 198850 389243
rect 1066 387589 198850 388155
rect 1066 386501 198850 387067
rect 1066 385413 198850 385979
rect 1066 384325 198850 384891
rect 1066 383237 198850 383803
rect 1066 382149 198850 382715
rect 1066 381061 198850 381627
rect 1066 379973 198850 380539
rect 1066 378885 198850 379451
rect 1066 377797 198850 378363
rect 1066 376709 198850 377275
rect 1066 375621 198850 376187
rect 1066 374533 198850 375099
rect 1066 373445 198850 374011
rect 1066 372357 198850 372923
rect 1066 371269 198850 371835
rect 1066 370181 198850 370747
rect 1066 369093 198850 369659
rect 1066 368005 198850 368571
rect 1066 366917 198850 367483
rect 1066 365829 198850 366395
rect 1066 364741 198850 365307
rect 1066 363653 198850 364219
rect 1066 362565 198850 363131
rect 1066 361477 198850 362043
rect 1066 360389 198850 360955
rect 1066 359301 198850 359867
rect 1066 358213 198850 358779
rect 1066 357125 198850 357691
rect 1066 356037 198850 356603
rect 1066 354949 198850 355515
rect 1066 353861 198850 354427
rect 1066 352773 198850 353339
rect 1066 351685 198850 352251
rect 1066 350597 198850 351163
rect 1066 349509 198850 350075
rect 1066 348421 198850 348987
rect 1066 347333 198850 347899
rect 1066 346245 198850 346811
rect 1066 345157 198850 345723
rect 1066 344069 198850 344635
rect 1066 342981 198850 343547
rect 1066 341893 198850 342459
rect 1066 340805 198850 341371
rect 1066 339717 198850 340283
rect 1066 338629 198850 339195
rect 1066 337541 198850 338107
rect 1066 336453 198850 337019
rect 1066 335365 198850 335931
rect 1066 334277 198850 334843
rect 1066 333189 198850 333755
rect 1066 332101 198850 332667
rect 1066 331013 198850 331579
rect 1066 329925 198850 330491
rect 1066 328837 198850 329403
rect 1066 327749 198850 328315
rect 1066 326661 198850 327227
rect 1066 325573 198850 326139
rect 1066 324485 198850 325051
rect 1066 323397 198850 323963
rect 1066 322309 198850 322875
rect 1066 321221 198850 321787
rect 1066 320133 198850 320699
rect 1066 319045 198850 319611
rect 1066 317957 198850 318523
rect 1066 316869 198850 317435
rect 1066 315781 198850 316347
rect 1066 314693 198850 315259
rect 1066 313605 198850 314171
rect 1066 312517 198850 313083
rect 1066 311429 198850 311995
rect 1066 310341 198850 310907
rect 1066 309253 198850 309819
rect 1066 308165 198850 308731
rect 1066 307077 198850 307643
rect 1066 305989 198850 306555
rect 1066 304901 198850 305467
rect 1066 303813 198850 304379
rect 1066 302725 198850 303291
rect 1066 301637 198850 302203
rect 1066 300549 198850 301115
rect 1066 299461 198850 300027
rect 1066 298373 198850 298939
rect 1066 297285 198850 297851
rect 1066 296197 198850 296763
rect 1066 295109 198850 295675
rect 1066 294021 198850 294587
rect 1066 292933 198850 293499
rect 1066 291845 198850 292411
rect 1066 290757 198850 291323
rect 1066 289669 198850 290235
rect 1066 288581 198850 289147
rect 1066 287493 198850 288059
rect 1066 286405 198850 286971
rect 1066 285317 198850 285883
rect 1066 284229 198850 284795
rect 1066 283141 198850 283707
rect 1066 282053 198850 282619
rect 1066 280965 198850 281531
rect 1066 279877 198850 280443
rect 1066 278789 198850 279355
rect 1066 277701 198850 278267
rect 1066 276613 198850 277179
rect 1066 275525 198850 276091
rect 1066 274437 198850 275003
rect 1066 273349 198850 273915
rect 1066 272261 198850 272827
rect 1066 271173 198850 271739
rect 1066 270085 198850 270651
rect 1066 268997 198850 269563
rect 1066 267909 198850 268475
rect 1066 266821 198850 267387
rect 1066 265733 198850 266299
rect 1066 264645 198850 265211
rect 1066 263557 198850 264123
rect 1066 262469 198850 263035
rect 1066 261381 198850 261947
rect 1066 260293 198850 260859
rect 1066 259205 198850 259771
rect 1066 258117 198850 258683
rect 1066 257029 198850 257595
rect 1066 255941 198850 256507
rect 1066 254853 198850 255419
rect 1066 253765 198850 254331
rect 1066 252677 198850 253243
rect 1066 251589 198850 252155
rect 1066 250501 198850 251067
rect 1066 249413 198850 249979
rect 1066 248325 198850 248891
rect 1066 247237 198850 247803
rect 1066 246149 198850 246715
rect 1066 245061 198850 245627
rect 1066 243973 198850 244539
rect 1066 242885 198850 243451
rect 1066 241797 198850 242363
rect 1066 240709 198850 241275
rect 1066 239621 198850 240187
rect 1066 238533 198850 239099
rect 1066 237445 198850 238011
rect 1066 236357 198850 236923
rect 1066 235269 198850 235835
rect 1066 234181 198850 234747
rect 1066 233093 198850 233659
rect 1066 232005 198850 232571
rect 1066 230917 198850 231483
rect 1066 229829 198850 230395
rect 1066 228741 198850 229307
rect 1066 227653 198850 228219
rect 1066 226565 198850 227131
rect 1066 225477 198850 226043
rect 1066 224389 198850 224955
rect 1066 223301 198850 223867
rect 1066 222213 198850 222779
rect 1066 221125 198850 221691
rect 1066 220037 198850 220603
rect 1066 218949 198850 219515
rect 1066 217861 198850 218427
rect 1066 216773 198850 217339
rect 1066 215685 198850 216251
rect 1066 214597 198850 215163
rect 1066 213509 198850 214075
rect 1066 212421 198850 212987
rect 1066 211333 198850 211899
rect 1066 210245 198850 210811
rect 1066 209157 198850 209723
rect 1066 208069 198850 208635
rect 1066 206981 198850 207547
rect 1066 205893 198850 206459
rect 1066 204805 198850 205371
rect 1066 203717 198850 204283
rect 1066 202629 198850 203195
rect 1066 201541 198850 202107
rect 1066 200453 198850 201019
rect 1066 199365 198850 199931
rect 1066 198277 198850 198843
rect 1066 197189 198850 197755
rect 1066 196101 198850 196667
rect 1066 195013 198850 195579
rect 1066 193925 198850 194491
rect 1066 192837 198850 193403
rect 1066 191749 198850 192315
rect 1066 190661 198850 191227
rect 1066 189573 198850 190139
rect 1066 188485 198850 189051
rect 1066 187397 198850 187963
rect 1066 186309 198850 186875
rect 1066 185221 198850 185787
rect 1066 184133 198850 184699
rect 1066 183045 198850 183611
rect 1066 181957 198850 182523
rect 1066 180869 198850 181435
rect 1066 179781 198850 180347
rect 1066 178693 198850 179259
rect 1066 177605 198850 178171
rect 1066 176517 198850 177083
rect 1066 175429 198850 175995
rect 1066 174341 198850 174907
rect 1066 173253 198850 173819
rect 1066 172165 198850 172731
rect 1066 171077 198850 171643
rect 1066 169989 198850 170555
rect 1066 168901 198850 169467
rect 1066 167813 198850 168379
rect 1066 166725 198850 167291
rect 1066 165637 198850 166203
rect 1066 164549 198850 165115
rect 1066 163461 198850 164027
rect 1066 162373 198850 162939
rect 1066 161285 198850 161851
rect 1066 160197 198850 160763
rect 1066 159109 198850 159675
rect 1066 158021 198850 158587
rect 1066 156933 198850 157499
rect 1066 155845 198850 156411
rect 1066 154757 198850 155323
rect 1066 153669 198850 154235
rect 1066 152581 198850 153147
rect 1066 151493 198850 152059
rect 1066 150405 198850 150971
rect 1066 149317 198850 149883
rect 1066 148229 198850 148795
rect 1066 147141 198850 147707
rect 1066 146053 198850 146619
rect 1066 144965 198850 145531
rect 1066 143877 198850 144443
rect 1066 142789 198850 143355
rect 1066 141701 198850 142267
rect 1066 140613 198850 141179
rect 1066 139525 198850 140091
rect 1066 138437 198850 139003
rect 1066 137349 198850 137915
rect 1066 136261 198850 136827
rect 1066 135173 198850 135739
rect 1066 134085 198850 134651
rect 1066 132997 198850 133563
rect 1066 131909 198850 132475
rect 1066 130821 198850 131387
rect 1066 129733 198850 130299
rect 1066 128645 198850 129211
rect 1066 127557 198850 128123
rect 1066 126469 198850 127035
rect 1066 125381 198850 125947
rect 1066 124293 198850 124859
rect 1066 123205 198850 123771
rect 1066 122117 198850 122683
rect 1066 121029 198850 121595
rect 1066 119941 198850 120507
rect 1066 118853 198850 119419
rect 1066 117765 198850 118331
rect 1066 116677 198850 117243
rect 1066 115589 198850 116155
rect 1066 114501 198850 115067
rect 1066 113413 198850 113979
rect 1066 112325 198850 112891
rect 1066 111237 198850 111803
rect 1066 110149 198850 110715
rect 1066 109061 198850 109627
rect 1066 107973 198850 108539
rect 1066 106885 198850 107451
rect 1066 105797 198850 106363
rect 1066 104709 198850 105275
rect 1066 103621 198850 104187
rect 1066 102533 198850 103099
rect 1066 101445 198850 102011
rect 1066 100357 198850 100923
rect 1066 99269 198850 99835
rect 1066 98181 198850 98747
rect 1066 97093 198850 97659
rect 1066 96005 198850 96571
rect 1066 94917 198850 95483
rect 1066 93829 198850 94395
rect 1066 92741 198850 93307
rect 1066 91653 198850 92219
rect 1066 90565 198850 91131
rect 1066 89477 198850 90043
rect 1066 88389 198850 88955
rect 1066 87301 198850 87867
rect 1066 86213 198850 86779
rect 1066 85125 198850 85691
rect 1066 84037 198850 84603
rect 1066 82949 198850 83515
rect 1066 81861 198850 82427
rect 1066 80773 198850 81339
rect 1066 79685 198850 80251
rect 1066 78597 198850 79163
rect 1066 77509 198850 78075
rect 1066 76421 198850 76987
rect 1066 75333 198850 75899
rect 1066 74245 198850 74811
rect 1066 73157 198850 73723
rect 1066 72069 198850 72635
rect 1066 70981 198850 71547
rect 1066 69893 198850 70459
rect 1066 68805 198850 69371
rect 1066 67717 198850 68283
rect 1066 66629 198850 67195
rect 1066 65541 198850 66107
rect 1066 64453 198850 65019
rect 1066 63365 198850 63931
rect 1066 62277 198850 62843
rect 1066 61189 198850 61755
rect 1066 60101 198850 60667
rect 1066 59013 198850 59579
rect 1066 57925 198850 58491
rect 1066 56837 198850 57403
rect 1066 55749 198850 56315
rect 1066 54661 198850 55227
rect 1066 53573 198850 54139
rect 1066 52485 198850 53051
rect 1066 51397 198850 51963
rect 1066 50309 198850 50875
rect 1066 49221 198850 49787
rect 1066 48133 198850 48699
rect 1066 47045 198850 47611
rect 1066 45957 198850 46523
rect 1066 44869 198850 45435
rect 1066 43781 198850 44347
rect 1066 42693 198850 43259
rect 1066 41605 198850 42171
rect 1066 40517 198850 41083
rect 1066 39429 198850 39995
rect 1066 38341 198850 38907
rect 1066 37253 198850 37819
rect 1066 36165 198850 36731
rect 1066 35077 198850 35643
rect 1066 33989 198850 34555
rect 1066 32901 198850 33467
rect 1066 31813 198850 32379
rect 1066 30725 198850 31291
rect 1066 29637 198850 30203
rect 1066 28549 198850 29115
rect 1066 27461 198850 28027
rect 1066 26373 198850 26939
rect 1066 25285 198850 25851
rect 1066 24197 198850 24763
rect 1066 23109 198850 23675
rect 1066 22021 198850 22587
rect 1066 20933 198850 21499
rect 1066 19845 198850 20411
rect 1066 18757 198850 19323
rect 1066 17669 198850 18235
rect 1066 16581 198850 17147
rect 1066 15493 198850 16059
rect 1066 14405 198850 14971
rect 1066 13317 198850 13883
rect 1066 12229 198850 12795
rect 1066 11141 198850 11707
rect 1066 10053 198850 10619
rect 1066 8965 198850 9531
rect 1066 7877 198850 8443
rect 1066 6789 198850 7355
rect 1066 5701 198850 6267
rect 1066 4613 198850 5179
rect 1066 3525 198850 4091
rect 1066 2437 198850 3003
<< obsli1 >>
rect 1104 2159 198812 397681
<< obsm1 >>
rect 1104 2048 198812 397712
<< metal2 >>
rect 49974 399200 50030 400000
rect 149978 399200 150034 400000
rect 2870 0 2926 800
rect 8574 0 8630 800
rect 14278 0 14334 800
rect 19982 0 20038 800
rect 25686 0 25742 800
rect 31390 0 31446 800
rect 37094 0 37150 800
rect 42798 0 42854 800
rect 48502 0 48558 800
rect 54298 0 54354 800
rect 60002 0 60058 800
rect 65706 0 65762 800
rect 71410 0 71466 800
rect 77114 0 77170 800
rect 82818 0 82874 800
rect 88522 0 88578 800
rect 94226 0 94282 800
rect 99930 0 99986 800
rect 105726 0 105782 800
rect 111430 0 111486 800
rect 117134 0 117190 800
rect 122838 0 122894 800
rect 128542 0 128598 800
rect 134246 0 134302 800
rect 139950 0 140006 800
rect 145654 0 145710 800
rect 151358 0 151414 800
rect 157154 0 157210 800
rect 162858 0 162914 800
rect 168562 0 168618 800
rect 174266 0 174322 800
rect 179970 0 180026 800
rect 185674 0 185730 800
rect 191378 0 191434 800
rect 197082 0 197138 800
<< obsm2 >>
rect 2872 399144 49918 399200
rect 50086 399144 149922 399200
rect 150090 399144 197964 399200
rect 2872 856 197964 399144
rect 2982 734 8518 856
rect 8686 734 14222 856
rect 14390 734 19926 856
rect 20094 734 25630 856
rect 25798 734 31334 856
rect 31502 734 37038 856
rect 37206 734 42742 856
rect 42910 734 48446 856
rect 48614 734 54242 856
rect 54410 734 59946 856
rect 60114 734 65650 856
rect 65818 734 71354 856
rect 71522 734 77058 856
rect 77226 734 82762 856
rect 82930 734 88466 856
rect 88634 734 94170 856
rect 94338 734 99874 856
rect 100042 734 105670 856
rect 105838 734 111374 856
rect 111542 734 117078 856
rect 117246 734 122782 856
rect 122950 734 128486 856
rect 128654 734 134190 856
rect 134358 734 139894 856
rect 140062 734 145598 856
rect 145766 734 151302 856
rect 151470 734 157098 856
rect 157266 734 162802 856
rect 162970 734 168506 856
rect 168674 734 174210 856
rect 174378 734 179914 856
rect 180082 734 185618 856
rect 185786 734 191322 856
rect 191490 734 197026 856
rect 197194 734 197964 856
<< obsm3 >>
rect 4208 2143 188848 397697
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
<< obsm4 >>
rect 34283 3435 34848 394093
rect 35328 3435 50208 394093
rect 50688 3435 65568 394093
rect 66048 3435 80928 394093
rect 81408 3435 96288 394093
rect 96768 3435 111648 394093
rect 112128 3435 127008 394093
rect 127488 3435 142368 394093
rect 142848 3435 157728 394093
rect 158208 3435 173088 394093
rect 173568 3435 173637 394093
<< labels >>
rlabel metal2 s 122838 0 122894 800 6 clk_i
port 1 nsew signal input
rlabel metal2 s 149978 399200 150034 400000 6 ds_n_o
port 2 nsew signal output
rlabel metal2 s 49974 399200 50030 400000 6 ds_o
port 3 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 fifo_ack_o
port 4 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 fifo_empty_o
port 5 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 fifo_full_o
port 6 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 fifo_i[0]
port 7 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 fifo_i[10]
port 8 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 fifo_i[11]
port 9 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 fifo_i[12]
port 10 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 fifo_i[13]
port 11 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 fifo_i[14]
port 12 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 fifo_i[15]
port 13 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 fifo_i[1]
port 14 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 fifo_i[2]
port 15 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 fifo_i[3]
port 16 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 fifo_i[4]
port 17 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 fifo_i[5]
port 18 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 fifo_i[6]
port 19 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 fifo_i[7]
port 20 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 fifo_i[8]
port 21 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 fifo_i[9]
port 22 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 fifo_rdy_i
port 23 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 mode_i
port 24 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 osr_i[0]
port 25 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 osr_i[1]
port 26 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 rst_n_i
port 27 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 tst_fifo_loop_i
port 28 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 tst_sinegen_en_i
port 29 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 tst_sinegen_step_i[0]
port 30 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 tst_sinegen_step_i[1]
port 31 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 tst_sinegen_step_i[2]
port 32 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 tst_sinegen_step_i[3]
port 33 nsew signal input
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 34 nsew power input
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 34 nsew power input
rlabel metal2 s 134246 0 134302 800 6 volume_i[0]
port 35 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 volume_i[1]
port 36 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 volume_i[2]
port 37 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 volume_i[3]
port 38 nsew signal input
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 39 nsew ground input
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 39 nsew ground input
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 39 nsew ground input
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 39 nsew ground input
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 39 nsew ground input
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 39 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 400000
string LEFview TRUE
string GDS_FILE /home/harald/caravel_mpw5/iic-audiodac-v1/openlane/audiodac/runs/audiodac/results/magic/audiodac.gds
string GDS_END 121227248
string GDS_START 697396
<< end >>

