`default_nettype none

module jku_logo(
	input jku
);

/* verilator lint_off UNUSED */
wire dummy1 = jku;
/* verilator lint_off UNUSED */

endmodule
`default_nettype wire
