VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO jku_logo
  CLASS BLOCK ;
  FOREIGN jku_logo ;
  ORIGIN -1.690 0.000 ;
  SIZE 1170.880 BY 376.070 ;
  PIN jku
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 541.715 90.355 545.140 90.360 ;
        RECT 344.570 5.505 747.425 90.355 ;
    END
  END jku
  OBS
      LAYER met4 ;
        RECT 186.855 147.495 272.570 376.070 ;
        RECT 344.570 369.140 346.285 372.605 ;
        RECT 744.780 371.250 747.425 372.605 ;
        RECT 344.570 367.410 349.715 369.140 ;
        RECT 744.000 367.410 747.425 371.250 ;
        RECT 344.570 363.950 354.855 367.410 ;
        RECT 742.285 365.680 747.425 367.410 ;
        RECT 738.855 363.950 747.425 365.680 ;
        RECT 344.570 362.215 353.140 363.950 ;
        RECT 735.425 362.215 747.425 363.950 ;
        RECT 344.570 360.485 356.570 362.215 ;
        RECT 733.715 360.485 747.425 362.215 ;
        RECT 344.570 358.755 358.285 360.485 ;
        RECT 732.000 358.755 747.425 360.485 ;
        RECT 344.570 357.020 361.715 358.755 ;
        RECT 730.285 357.020 747.425 358.755 ;
        RECT 344.570 353.560 366.855 357.020 ;
        RECT 728.570 355.290 747.425 357.020 ;
        RECT 726.855 353.560 747.425 355.290 ;
        RECT 344.570 351.825 368.570 353.560 ;
        RECT 723.425 351.825 747.425 353.560 ;
        RECT 344.570 350.095 370.285 351.825 ;
        RECT 720.000 350.095 747.425 351.825 ;
        RECT 344.570 348.365 372.000 350.095 ;
        RECT 721.715 348.365 747.425 350.095 ;
        RECT 344.570 346.630 373.715 348.365 ;
        RECT 344.570 344.900 377.140 346.630 ;
        RECT 718.285 344.900 747.425 348.365 ;
        RECT 344.570 341.435 378.855 344.900 ;
        RECT 714.855 343.170 747.425 344.900 ;
        RECT 713.140 341.435 747.425 343.170 ;
        RECT 344.570 337.975 382.285 341.435 ;
        RECT 709.715 339.705 747.425 341.435 ;
        RECT 708.000 337.975 747.425 339.705 ;
        RECT 344.570 336.240 385.715 337.975 ;
        RECT 706.285 336.240 747.425 337.975 ;
        RECT 344.570 334.510 387.425 336.240 ;
        RECT 704.570 334.510 747.425 336.240 ;
        RECT 344.570 332.780 390.855 334.510 ;
        RECT 702.855 332.780 747.425 334.510 ;
        RECT 344.570 331.045 392.570 332.780 ;
        RECT 699.425 331.045 747.425 332.780 ;
        RECT 344.570 329.315 394.285 331.045 ;
        RECT 696.000 329.315 747.425 331.045 ;
        RECT 344.570 327.585 396.000 329.315 ;
        RECT 697.715 327.585 747.425 329.315 ;
        RECT 344.570 325.850 397.715 327.585 ;
        RECT 344.570 324.120 401.140 325.850 ;
        RECT 694.285 324.120 747.425 327.585 ;
        RECT 344.570 320.660 402.855 324.120 ;
        RECT 692.570 322.390 747.425 324.120 ;
        RECT 689.140 320.660 747.425 322.390 ;
        RECT 344.570 318.925 404.570 320.660 ;
        RECT 685.715 318.925 747.425 320.660 ;
        RECT 344.570 317.195 406.285 318.925 ;
        RECT 684.000 317.195 747.425 318.925 ;
        RECT 344.570 315.465 408.000 317.195 ;
        RECT 682.285 315.465 747.425 317.195 ;
        RECT 344.570 313.730 411.425 315.465 ;
        RECT 413.140 313.730 414.855 315.465 ;
        RECT 344.570 312.000 414.855 313.730 ;
        RECT 677.140 312.000 678.855 313.730 ;
        RECT 680.570 312.000 747.425 315.465 ;
        RECT 344.570 310.270 416.570 312.000 ;
        RECT 677.140 310.270 747.425 312.000 ;
        RECT 344.570 308.535 418.285 310.270 ;
        RECT 673.715 308.535 747.425 310.270 ;
        RECT 344.570 305.075 420.000 308.535 ;
        RECT 421.715 305.075 423.425 306.805 ;
        RECT 672.000 305.075 747.425 308.535 ;
        RECT 344.570 301.610 425.140 305.075 ;
        RECT 668.570 301.610 747.425 305.075 ;
        RECT 344.570 298.145 428.570 301.610 ;
        RECT 665.140 299.880 747.425 301.610 ;
        RECT 344.570 294.685 432.000 298.145 ;
        RECT 660.000 296.415 747.425 299.880 ;
        RECT 433.715 294.685 435.425 296.415 ;
        RECT 658.285 294.685 747.425 296.415 ;
        RECT 344.570 291.220 438.855 294.685 ;
        RECT 656.570 292.950 747.425 294.685 ;
        RECT 654.855 291.220 747.425 292.950 ;
        RECT 344.570 289.490 440.570 291.220 ;
        RECT 653.140 289.490 747.425 291.220 ;
        RECT 344.570 287.755 442.285 289.490 ;
        RECT 648.000 287.755 649.715 289.490 ;
        RECT 651.425 287.755 747.425 289.490 ;
        RECT 344.570 286.025 444.000 287.755 ;
        RECT 344.570 284.295 447.425 286.025 ;
        RECT 648.000 284.295 747.425 287.755 ;
        RECT 344.570 280.830 449.140 284.295 ;
        RECT 641.140 280.830 642.855 282.560 ;
        RECT 644.570 280.830 747.425 284.295 ;
        RECT 344.570 277.365 452.570 280.830 ;
        RECT 641.140 279.100 747.425 280.830 ;
        RECT 344.570 275.635 454.285 277.365 ;
        RECT 636.000 275.635 747.425 279.100 ;
        RECT 344.570 273.905 456.000 275.635 ;
        RECT 457.715 273.905 459.425 275.635 ;
        RECT 634.285 273.905 747.425 275.635 ;
        RECT 344.570 270.440 462.855 273.905 ;
        RECT 632.570 272.175 747.425 273.905 ;
        RECT 630.855 270.440 747.425 272.175 ;
        RECT 346.285 268.710 464.570 270.440 ;
        RECT 629.140 268.710 747.425 270.440 ;
        RECT 348.000 266.980 466.285 268.710 ;
        RECT 624.000 266.980 744.000 268.710 ;
        RECT 349.715 265.245 468.000 266.980 ;
        RECT 624.000 265.280 740.930 266.980 ;
        RECT 624.000 265.245 738.855 265.280 ;
        RECT 351.425 263.515 469.715 265.245 ;
        RECT 622.285 263.515 738.855 265.245 ;
        RECT 353.140 261.785 473.140 263.515 ;
        RECT 622.285 261.785 737.140 263.515 ;
        RECT 356.570 260.050 476.570 261.785 ;
        RECT 620.570 260.790 735.425 261.785 ;
        RECT 620.570 260.050 735.410 260.790 ;
        RECT 358.285 258.320 474.855 260.050 ;
        RECT 615.425 258.320 617.140 260.050 ;
        RECT 618.855 258.320 735.410 260.050 ;
        RECT 361.715 254.855 478.285 258.320 ;
        RECT 615.425 256.590 733.715 258.320 ;
        RECT 612.000 254.855 730.285 256.590 ;
        RECT 361.715 253.125 363.425 254.855 ;
        RECT 365.140 253.410 483.425 254.855 ;
        RECT 365.140 253.125 483.430 253.410 ;
        RECT 610.285 253.125 728.570 254.855 ;
        RECT 365.140 251.395 485.140 253.125 ;
        RECT 608.570 251.395 726.855 253.125 ;
        RECT 366.855 249.660 486.855 251.395 ;
        RECT 606.855 249.660 725.140 251.395 ;
        RECT 370.285 247.930 488.570 249.660 ;
        RECT 605.140 247.930 723.425 249.660 ;
        RECT 372.000 246.200 490.285 247.930 ;
        RECT 600.000 246.200 720.000 247.930 ;
        RECT 373.715 244.465 492.000 246.200 ;
        RECT 601.715 244.465 718.285 246.200 ;
        RECT 375.425 242.735 493.715 244.465 ;
        RECT 375.425 241.005 377.140 242.735 ;
        RECT 378.855 241.005 497.140 242.735 ;
        RECT 598.285 241.005 714.855 244.465 ;
        RECT 380.570 239.270 498.855 241.005 ;
        RECT 593.140 240.070 711.425 241.005 ;
        RECT 593.140 239.270 711.190 240.070 ;
        RECT 382.285 237.540 498.855 239.270 ;
        RECT 594.855 237.540 711.190 239.270 ;
        RECT 385.715 234.075 502.285 237.540 ;
        RECT 589.715 235.810 709.715 237.540 ;
        RECT 588.000 234.075 706.285 235.810 ;
        RECT 387.425 232.350 507.425 234.075 ;
        RECT 387.425 232.345 507.430 232.350 ;
        RECT 586.285 232.345 704.570 234.075 ;
        RECT 389.140 230.615 509.140 232.345 ;
        RECT 584.570 230.615 702.855 232.345 ;
        RECT 390.855 228.885 510.855 230.615 ;
        RECT 582.855 228.885 701.140 230.615 ;
        RECT 394.285 227.150 512.570 228.885 ;
        RECT 579.425 227.150 697.715 228.885 ;
        RECT 396.000 225.420 514.285 227.150 ;
        RECT 577.715 225.420 696.000 227.150 ;
        RECT 397.715 223.690 516.000 225.420 ;
        RECT 576.000 223.690 694.285 225.420 ;
        RECT 399.425 221.955 517.715 223.690 ;
        RECT 574.285 222.550 691.550 223.690 ;
        RECT 399.425 221.910 401.140 221.955 ;
        RECT 402.855 220.225 521.140 221.955 ;
        RECT 574.285 220.225 689.140 222.550 ;
        RECT 404.570 218.495 522.855 220.225 ;
        RECT 572.570 218.495 687.060 220.225 ;
        RECT 406.285 216.760 522.855 218.495 ;
        RECT 569.140 218.160 687.060 218.495 ;
        RECT 409.715 215.030 526.285 216.760 ;
        RECT 565.715 215.030 567.425 216.760 ;
        RECT 569.140 215.030 685.715 218.160 ;
        RECT 411.425 213.300 526.285 215.030 ;
        RECT 564.000 213.300 682.285 215.030 ;
        RECT 411.425 211.565 529.715 213.300 ;
        RECT 562.285 211.565 680.570 213.300 ;
        RECT 412.760 211.100 533.140 211.565 ;
        RECT 413.140 209.835 533.140 211.100 ;
        RECT 560.570 209.835 678.855 211.565 ;
        RECT 414.855 208.105 416.570 209.835 ;
        RECT 418.285 208.105 534.855 209.835 ;
        RECT 558.855 208.105 677.140 209.835 ;
        RECT 418.285 206.370 536.570 208.105 ;
        RECT 557.140 206.370 673.715 208.105 ;
        RECT 421.715 204.640 538.285 206.370 ;
        RECT 552.000 204.640 672.000 206.370 ;
        RECT 421.715 202.910 540.000 204.640 ;
        RECT 552.000 202.910 670.285 204.640 ;
        RECT 423.425 201.175 543.425 202.910 ;
        RECT 552.000 201.175 666.855 202.910 ;
        RECT 426.855 199.445 545.140 201.175 ;
        RECT 548.570 199.445 665.140 201.175 ;
        RECT 428.570 197.715 665.140 199.445 ;
        RECT 430.285 195.980 661.715 197.715 ;
        RECT 663.425 197.650 665.140 197.715 ;
        RECT 432.000 194.250 661.715 195.980 ;
        RECT 435.425 192.520 660.000 194.250 ;
        RECT 437.140 190.785 656.570 192.520 ;
        RECT 438.855 189.055 654.855 190.785 ;
        RECT 440.570 187.240 653.140 189.055 ;
        RECT 440.570 185.595 651.700 187.240 ;
        RECT 444.000 183.860 648.000 185.595 ;
        RECT 445.715 182.130 646.285 183.860 ;
        RECT 819.425 182.130 903.425 376.070 ;
        RECT 447.425 180.400 644.570 182.130 ;
        RECT 449.140 178.665 641.140 180.400 ;
        RECT 452.570 176.935 641.140 178.665 ;
        RECT 819.425 176.935 905.140 182.130 ;
        RECT 454.285 175.205 641.140 176.935 ;
        RECT 821.140 175.205 905.140 176.935 ;
        RECT 1086.855 178.665 1170.855 376.070 ;
        RECT 1086.855 175.205 1172.570 178.665 ;
        RECT 456.000 173.470 637.715 175.205 ;
        RECT 459.425 171.770 636.000 173.470 ;
        RECT 459.425 170.010 632.570 171.770 ;
        RECT 634.285 171.740 636.000 171.770 ;
        RECT 819.425 171.740 906.855 175.205 ;
        RECT 464.570 168.275 630.855 170.010 ;
        RECT 819.425 168.275 905.140 171.740 ;
        RECT 1086.855 170.010 1170.855 175.205 ;
        RECT 462.855 166.545 629.140 168.275 ;
        RECT 468.000 164.815 627.425 166.545 ;
        RECT 468.000 163.080 624.000 164.815 ;
        RECT 471.425 161.350 622.285 163.080 ;
        RECT 821.140 161.350 905.140 168.275 ;
        RECT 1085.140 166.545 1170.855 170.010 ;
        RECT 1085.140 164.815 1169.140 166.545 ;
        RECT 1083.425 163.080 1169.140 164.815 ;
        RECT 471.425 159.620 620.570 161.350 ;
        RECT 471.425 157.885 615.425 159.620 ;
        RECT 476.570 156.155 615.425 157.885 ;
        RECT 478.285 154.425 615.520 156.155 ;
        RECT 480.000 153.680 613.920 154.425 ;
        RECT 480.000 152.690 613.715 153.680 ;
        RECT 485.140 149.230 608.570 152.690 ;
        RECT 821.140 149.230 906.855 161.350 ;
        RECT 1085.140 152.690 1169.140 163.080 ;
        RECT 1081.715 150.960 1169.140 152.690 ;
        RECT 1083.425 149.230 1170.855 150.960 ;
        RECT 485.140 147.495 605.140 149.230 ;
        RECT 821.140 147.495 908.570 149.230 ;
        RECT 185.140 131.915 272.570 147.495 ;
        RECT 486.855 145.765 605.140 147.495 ;
        RECT 490.285 144.035 603.425 145.765 ;
        RECT 492.000 142.305 600.000 144.035 ;
        RECT 493.715 140.570 598.285 142.305 ;
        RECT 822.855 140.570 908.570 147.495 ;
        RECT 1083.425 147.495 1169.140 149.230 ;
        RECT 1083.425 145.765 1167.425 147.495 ;
        RECT 495.425 138.840 596.570 140.570 ;
        RECT 495.425 137.110 594.855 138.840 ;
        RECT 500.570 135.375 593.280 137.110 ;
        RECT 502.285 134.470 593.280 135.375 ;
        RECT 822.855 135.375 910.285 140.570 ;
        RECT 1081.715 138.840 1167.425 145.765 ;
        RECT 1080.000 137.110 1169.140 138.840 ;
        RECT 1080.000 135.375 1167.425 137.110 ;
        RECT 502.285 133.645 593.140 134.470 ;
        RECT 822.855 133.645 912.000 135.375 ;
        RECT 1080.000 133.645 1165.715 135.375 ;
        RECT 185.140 130.180 272.600 131.915 ;
        RECT 505.715 130.180 586.285 133.645 ;
        RECT 588.000 131.915 589.715 133.645 ;
        RECT 824.570 131.915 912.000 133.645 ;
        RECT 1078.285 131.915 1165.715 133.645 ;
        RECT 183.425 126.720 272.570 130.180 ;
        RECT 509.140 126.720 582.855 130.180 ;
        RECT 824.570 126.720 913.715 131.915 ;
        RECT 1080.000 130.180 1165.715 131.915 ;
        RECT 1078.285 128.450 1165.715 130.180 ;
        RECT 183.425 121.525 270.855 126.720 ;
        RECT 510.855 124.985 581.140 126.720 ;
        RECT 826.285 124.985 915.425 126.720 ;
        RECT 1076.570 124.985 1165.715 128.450 ;
        RECT 514.285 123.255 579.425 124.985 ;
        RECT 516.000 121.525 577.715 123.255 ;
        RECT 826.285 121.525 917.140 124.985 ;
        RECT 1074.855 121.525 1164.000 124.985 ;
        RECT 53.140 118.060 54.855 119.790 ;
        RECT 51.425 116.330 58.285 118.060 ;
        RECT 181.715 116.330 270.855 121.525 ;
        RECT 517.715 119.790 574.285 121.525 ;
        RECT 521.140 118.060 572.570 119.790 ;
        RECT 826.285 118.060 918.855 121.525 ;
        RECT 1073.140 119.790 1164.000 121.525 ;
        RECT 1073.140 118.060 1162.285 119.790 ;
        RECT 522.855 116.330 570.855 118.060 ;
        RECT 49.715 114.610 60.000 116.330 ;
        RECT 47.190 114.595 60.000 114.610 ;
        RECT 181.660 114.595 270.855 116.330 ;
        RECT 524.570 114.595 565.715 116.330 ;
        RECT 47.190 112.865 61.715 114.595 ;
        RECT 181.715 112.865 270.855 114.595 ;
        RECT 526.285 112.865 565.715 114.595 ;
        RECT 828.000 114.595 920.570 118.060 ;
        RECT 1071.425 116.330 1162.285 118.060 ;
        RECT 828.000 112.865 922.285 114.595 ;
        RECT 1069.715 112.865 1162.285 116.330 ;
        RECT 45.910 111.190 63.425 112.865 ;
        RECT 44.100 109.400 63.425 111.190 ;
        RECT 180.000 111.135 270.855 112.865 ;
        RECT 531.425 111.135 565.715 112.865 ;
        RECT 829.715 111.135 924.000 112.865 ;
        RECT 42.855 107.670 65.140 109.400 ;
        RECT 178.285 107.760 269.140 111.135 ;
        RECT 531.425 110.340 564.270 111.135 ;
        RECT 531.425 109.400 564.000 110.340 ;
        RECT 178.285 107.670 268.980 107.760 ;
        RECT 534.855 107.670 558.855 109.400 ;
        RECT 41.140 106.110 66.855 107.670 ;
        RECT 41.130 105.940 66.855 106.110 ;
        RECT 41.130 104.205 68.570 105.940 ;
        RECT 176.570 104.205 268.980 107.670 ;
        RECT 534.550 105.940 558.855 107.670 ;
        RECT 829.715 107.670 925.715 111.135 ;
        RECT 1068.000 109.400 1160.570 112.865 ;
        RECT 1064.570 107.670 1162.285 109.400 ;
        RECT 829.715 105.940 927.425 107.670 ;
        RECT 1062.855 105.940 1158.855 107.670 ;
        RECT 538.285 104.205 555.425 105.940 ;
        RECT 831.425 104.205 929.140 105.940 ;
        RECT 1064.570 104.205 1158.855 105.940 ;
        RECT 39.425 102.475 70.285 104.205 ;
        RECT 174.855 103.340 268.980 104.205 ;
        RECT 174.855 102.475 269.140 103.340 ;
        RECT 538.060 102.475 555.470 104.205 ;
        RECT 37.715 100.745 72.000 102.475 ;
        RECT 173.140 101.430 267.425 102.475 ;
        RECT 36.000 99.130 75.900 100.745 ;
        RECT 36.000 99.015 77.140 99.130 ;
        RECT 34.285 97.280 77.140 99.015 ;
        RECT 173.040 98.280 267.425 101.430 ;
        RECT 541.715 100.745 553.715 102.475 ;
        RECT 831.425 100.745 932.570 104.205 ;
        RECT 1061.140 102.475 1158.855 104.205 ;
        RECT 1061.140 100.745 1157.140 102.475 ;
        RECT 541.715 99.015 550.285 100.745 ;
        RECT 833.140 99.015 934.285 100.745 ;
        RECT 1056.000 99.015 1157.140 100.745 ;
        RECT 173.140 97.280 267.425 98.280 ;
        RECT 543.425 97.280 548.570 99.015 ;
        RECT 833.140 97.280 936.000 99.015 ;
        RECT 1057.715 97.280 1157.140 99.015 ;
        RECT 32.570 95.550 80.570 97.280 ;
        RECT 169.715 95.550 267.425 97.280 ;
        RECT 833.140 95.580 939.425 97.280 ;
        RECT 833.140 95.550 939.450 95.580 ;
        RECT 1052.570 95.550 1155.425 97.280 ;
        RECT 30.220 94.620 82.285 95.550 ;
        RECT 29.140 93.820 82.285 94.620 ;
        RECT 168.000 93.820 265.715 95.550 ;
        RECT 29.140 92.085 84.000 93.820 ;
        RECT 27.425 90.355 85.715 92.085 ;
        RECT 166.360 91.480 265.715 93.820 ;
        RECT 834.855 92.085 942.855 95.550 ;
        RECT 1054.285 93.820 1155.425 95.550 ;
        RECT 1049.140 92.085 1153.715 93.820 ;
        RECT 166.285 90.355 265.715 91.480 ;
        RECT 836.570 90.355 946.285 92.085 ;
        RECT 1045.715 90.355 1153.715 92.085 ;
        RECT 27.425 88.625 89.140 90.355 ;
        RECT 161.140 88.920 264.000 90.355 ;
        RECT 25.715 86.890 94.285 88.625 ;
        RECT 160.630 86.890 264.000 88.920 ;
        RECT 836.570 88.625 948.000 90.355 ;
        RECT 1044.000 88.625 1153.715 90.355 ;
        RECT 24.000 85.160 96.000 86.890 ;
        RECT 157.715 85.160 264.000 86.890 ;
        RECT 838.285 86.890 948.000 88.625 ;
        RECT 1038.855 86.890 1152.000 88.625 ;
        RECT 838.285 85.160 954.855 86.890 ;
        RECT 1037.140 85.160 1152.000 86.890 ;
        RECT 22.285 83.430 99.425 85.160 ;
        RECT 152.570 83.430 154.285 83.470 ;
        RECT 156.000 83.430 262.285 85.160 ;
        RECT 20.570 81.695 106.285 83.430 ;
        RECT 144.000 81.695 145.715 81.700 ;
        RECT 149.140 81.695 262.285 83.430 ;
        RECT 840.000 83.430 960.000 85.160 ;
        RECT 1032.000 83.430 1150.285 85.160 ;
        RECT 840.000 81.695 963.425 83.430 ;
        RECT 1026.855 81.695 1150.285 83.430 ;
        RECT 18.855 79.965 109.715 81.695 ;
        RECT 111.425 79.965 114.855 81.695 ;
        RECT 142.285 79.965 262.410 81.695 ;
        RECT 841.715 79.965 972.000 81.695 ;
        RECT 1020.000 79.965 1148.570 81.695 ;
        RECT 18.855 79.320 260.570 79.965 ;
        RECT 16.400 76.500 260.570 79.320 ;
        RECT 841.715 78.235 980.570 79.965 ;
        RECT 1011.425 78.235 1148.570 79.965 ;
        RECT 13.715 74.770 260.570 76.500 ;
        RECT 843.425 74.770 1146.855 78.235 ;
        RECT 15.425 73.040 258.855 74.770 ;
        RECT 12.000 71.305 258.855 73.040 ;
        RECT 845.140 71.305 1145.140 74.770 ;
        RECT 8.570 71.180 10.285 71.305 ;
        RECT 12.000 71.180 257.140 71.305 ;
        RECT 8.570 69.575 257.140 71.180 ;
        RECT 846.855 70.130 1145.140 71.305 ;
        RECT 846.855 69.575 1141.715 70.130 ;
        RECT 1143.425 69.575 1145.140 70.130 ;
        RECT 8.570 67.845 255.425 69.575 ;
        RECT 6.855 66.110 255.425 67.845 ;
        RECT 850.285 67.845 1141.715 69.575 ;
        RECT 850.285 66.110 1141.620 67.845 ;
        RECT 5.140 64.380 255.450 66.110 ;
        RECT 850.285 64.380 1141.715 66.110 ;
        RECT 3.425 62.650 253.715 64.380 ;
        RECT 1.715 60.915 253.715 62.650 ;
        RECT 852.000 60.915 1138.285 64.380 ;
        RECT 1.690 59.185 252.000 60.915 ;
        RECT 853.715 59.185 1136.570 60.915 ;
        RECT 3.425 57.455 250.285 59.185 ;
        RECT 5.140 55.720 250.285 57.455 ;
        RECT 855.425 57.455 1134.855 59.185 ;
        RECT 855.425 55.720 1133.140 57.455 ;
        RECT 5.140 53.990 248.570 55.720 ;
        RECT 855.425 53.990 857.140 55.720 ;
        RECT 858.855 53.990 1131.425 55.720 ;
        RECT 6.855 52.360 248.570 53.990 ;
        RECT 6.855 52.260 246.130 52.360 ;
        RECT 860.570 52.260 1129.715 53.990 ;
        RECT 8.570 50.530 245.140 52.260 ;
        RECT 10.285 48.795 245.140 50.530 ;
        RECT 864.000 50.530 1129.715 52.260 ;
        RECT 12.000 47.065 243.425 48.795 ;
        RECT 864.000 47.065 1128.000 50.530 ;
        RECT 13.715 45.335 241.715 47.065 ;
        RECT 865.715 45.335 1126.285 47.065 ;
        RECT 15.425 43.600 241.715 45.335 ;
        RECT 867.425 43.600 1124.570 45.335 ;
        RECT 17.140 41.870 240.000 43.600 ;
        RECT 869.140 41.870 1121.140 43.600 ;
        RECT 18.855 40.140 238.285 41.870 ;
        RECT 872.570 40.140 1119.425 41.870 ;
        RECT 19.830 40.100 236.570 40.140 ;
        RECT 22.285 38.405 236.570 40.100 ;
        RECT 874.285 38.405 1116.000 40.140 ;
        RECT 22.285 36.675 234.855 38.405 ;
        RECT 874.285 36.675 876.000 38.405 ;
        RECT 877.715 36.675 1114.285 38.405 ;
        RECT 25.715 34.945 233.140 36.675 ;
        RECT 874.285 34.945 1112.570 36.675 ;
        RECT 27.425 33.210 231.425 34.945 ;
        RECT 881.140 33.210 1110.855 34.945 ;
        RECT 29.140 31.480 229.715 33.210 ;
        RECT 881.140 31.480 1109.140 33.210 ;
        RECT 30.855 29.750 228.000 31.480 ;
        RECT 882.855 29.750 1105.715 31.480 ;
        RECT 31.600 29.610 226.285 29.750 ;
        RECT 36.000 28.230 226.285 29.610 ;
        RECT 36.000 26.285 222.855 28.230 ;
        RECT 224.570 28.015 226.285 28.230 ;
        RECT 886.285 28.015 1104.000 29.750 ;
        RECT 888.000 26.285 1100.570 28.015 ;
        RECT 39.425 24.555 222.855 26.285 ;
        RECT 891.425 24.555 1100.570 26.285 ;
        RECT 42.855 22.820 217.715 24.555 ;
        RECT 894.855 22.820 1095.425 24.555 ;
        RECT 46.285 21.090 214.285 22.820 ;
        RECT 898.285 21.090 1090.285 22.820 ;
        RECT 48.000 19.360 212.570 21.090 ;
        RECT 900.000 19.360 1088.570 21.090 ;
        RECT 53.140 17.625 209.140 19.360 ;
        RECT 905.140 17.625 1085.140 19.360 ;
        RECT 54.855 15.895 205.715 17.625 ;
        RECT 908.570 15.895 1081.715 17.625 ;
        RECT 58.285 14.165 202.285 15.895 ;
        RECT 910.285 14.165 1078.285 15.895 ;
        RECT 63.425 12.430 198.855 14.165 ;
        RECT 200.570 13.920 202.285 14.165 ;
        RECT 915.425 12.430 1073.140 14.165 ;
        RECT 66.855 10.700 192.000 12.430 ;
        RECT 193.715 12.250 195.425 12.430 ;
        RECT 920.570 10.700 1068.000 12.430 ;
        RECT 72.000 8.970 188.570 10.700 ;
        RECT 925.715 8.970 1062.855 10.700 ;
        RECT 1066.285 8.970 1068.000 10.700 ;
        RECT 77.140 7.240 185.140 8.970 ;
        RECT 930.855 7.240 932.570 8.970 ;
        RECT 934.285 7.240 1054.285 8.970 ;
        RECT 1056.000 7.240 1057.715 8.970 ;
        RECT 84.000 5.505 178.285 7.240 ;
        RECT 937.715 5.505 1050.855 7.240 ;
        RECT 90.855 3.775 171.425 5.505 ;
        RECT 944.570 3.775 946.285 5.505 ;
        RECT 948.000 3.775 1044.000 5.505 ;
        RECT 101.140 2.045 161.140 3.775 ;
        RECT 956.570 2.045 1032.000 3.775 ;
        RECT 102.855 1.860 104.570 2.045 ;
        RECT 114.855 0.310 147.425 2.045 ;
        RECT 157.715 1.960 159.425 2.045 ;
        RECT 966.855 0.310 1014.855 2.045 ;
        RECT 1016.570 0.310 1021.715 2.045 ;
        RECT 121.715 0.000 123.425 0.310 ;
        RECT 138.855 0.000 140.570 0.310 ;
  END
END jku_logo
END LIBRARY

